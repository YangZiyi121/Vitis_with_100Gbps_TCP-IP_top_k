   
    parameter PROC_NUM = 69;
    parameter ST_IDLE = 3'b000;
    parameter ST_FILTER_FAKE = 3'b001;
    parameter ST_DL_DETECTED = 3'b010;
    parameter ST_DL_REPORT = 3'b100;
   

    reg [2:0] CS_fsm;
    reg [2:0] NS_fsm;
    reg [PROC_NUM - 1:0] dl_detect_reg;
    reg [PROC_NUM - 1:0] dl_done_reg;
    reg [PROC_NUM - 1:0] origin_reg;
    reg [PROC_NUM - 1:0] dl_in_vec_reg;
    reg [31:0] dl_keep_cnt;
    integer i;
    integer fp;

    // FSM State machine
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            CS_fsm <= ST_IDLE;
        end
        else begin
            CS_fsm <= NS_fsm;
        end
    end
    always @ (CS_fsm or dl_in_vec or dl_detect_reg or dl_done_reg or dl_in_vec or origin_reg or dl_keep_cnt) begin
        case (CS_fsm)
            ST_IDLE : begin
                if (|dl_in_vec) begin
                    NS_fsm = ST_FILTER_FAKE;
                end
                else begin
                    NS_fsm = ST_IDLE;
                end
            end
            ST_FILTER_FAKE: begin
                if (dl_keep_cnt >= 32'd1000) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else if (dl_detect_reg != (dl_detect_reg & dl_in_vec)) begin
                    NS_fsm = ST_IDLE;
                end
                else begin
                    NS_fsm = ST_FILTER_FAKE;
                end
            end
            ST_DL_DETECTED: begin
                // has unreported deadlock cycle
                if (dl_detect_reg != dl_done_reg) begin
                    NS_fsm = ST_DL_REPORT;
                end
                else begin
                    NS_fsm = ST_DL_DETECTED;
                end
            end
            ST_DL_REPORT: begin
                if (|(dl_in_vec & origin_reg)) begin
                    NS_fsm = ST_DL_DETECTED;
                end
                else begin
                    NS_fsm = ST_DL_REPORT;
                end
            end
            default: NS_fsm = ST_IDLE;
        endcase
    end

    // dl_detect_reg record the procs that first detect deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_detect_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_IDLE) begin
                dl_detect_reg <= dl_in_vec;
            end
        end
    end

    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_keep_cnt <= 32'h0;
        end
        else begin
            if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg == (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= dl_keep_cnt + 32'h1;
            end
            else if (CS_fsm == ST_FILTER_FAKE && (dl_detect_reg != (dl_detect_reg & dl_in_vec))) begin
                dl_keep_cnt <= 32'h0;
            end
        end
    end

    // dl_detect_out keeps in high after deadlock detected
    assign dl_detect_out = (|dl_detect_reg) && (CS_fsm == ST_DL_DETECTED || CS_fsm == ST_DL_REPORT);

    // dl_done_reg record the cycles has been reported
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_done_reg <= 'b0;
        end
        else begin
            if ((CS_fsm == ST_DL_REPORT) && (|(dl_in_vec & dl_detect_reg) == 'b1)) begin
                dl_done_reg <= dl_done_reg | dl_in_vec;
            end
        end
    end

    // clear token once a cycle is done
    assign token_clear = (CS_fsm == ST_DL_REPORT) ? ((|(dl_in_vec & origin_reg)) ? 'b1 : 'b0) : 'b0;

    // origin_reg record the current cycle start id
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            origin_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                origin_reg <= origin;
            end
        end
    end
   
    // origin will be valid for only one cycle
    wire [PROC_NUM*PROC_NUM - 1:0] origin_tmp;
    assign origin_tmp[PROC_NUM - 1:0] = (dl_detect_reg[0] & ~dl_done_reg[0]) ? 'b1 : 'b0;
    genvar j;
    generate
    for(j = 1;j < PROC_NUM;j = j + 1) begin: F1
        assign origin_tmp[j*PROC_NUM +: PROC_NUM] = (dl_detect_reg[j] & ~dl_done_reg[j]) ? ('b1 << j) : origin_tmp[(j - 1)*PROC_NUM +: PROC_NUM];
    end
    endgenerate
    always @ (CS_fsm or origin_tmp) begin
        if (CS_fsm == ST_DL_DETECTED) begin
            origin = origin_tmp[(PROC_NUM - 1)*PROC_NUM +: PROC_NUM];
        end
        else begin
            origin = 'b0;
        end
    end

    
    // dl_in_vec_reg record the current cycle dl_in_vec
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            dl_in_vec_reg <= 'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED) begin
                dl_in_vec_reg <= origin;
            end
            else if (CS_fsm == ST_DL_REPORT) begin
                dl_in_vec_reg <= dl_in_vec;
            end
        end
    end
    
    // find_df_deadlock to report the deadlock
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            find_df_deadlock <= 1'b0;
        end
        else begin
            if (CS_fsm == ST_DL_DETECTED && dl_detect_reg == dl_done_reg) begin
                find_df_deadlock <= 1'b1;
            end
            else if (CS_fsm == ST_IDLE) begin
                find_df_deadlock <= 1'b0;
            end
        end
    end
    
    // get the first valid proc index in dl vector
    function integer proc_index(input [PROC_NUM - 1:0] dl_vec);
        begin
            proc_index = 0;
            for (i = 0; i < PROC_NUM; i = i + 1) begin
                if (dl_vec[i]) begin
                    proc_index = i;
                end
            end
        end
    endfunction

    // get the proc path based on dl vector
    function [488:0] proc_path(input [PROC_NUM - 1:0] dl_vec);
        integer index;
        begin
            index = proc_index(dl_vec);
            case (index)
                0 : begin
                    proc_path = "toe_top_toe_top.entry_proc_U0";
                end
                1 : begin
                    proc_path = "toe_top_toe_top.convert_axis_to_net_axis_512_U0";
                end
                2 : begin
                    proc_path = "toe_top_toe_top.convert_axis_to_net_axis_512_1_U0";
                end
                3 : begin
                    proc_path = "toe_top_toe_top.convert_axis_to_net_axis_512_2_U0";
                end
                4 : begin
                    proc_path = "toe_top_toe_top.convert_net_axis_to_axis_512_U0";
                end
                5 : begin
                    proc_path = "toe_top_toe_top.convert_net_axis_to_axis_512_1_U0";
                end
                6 : begin
                    proc_path = "toe_top_toe_top.convert_net_axis_to_axis_512_2_U0";
                end
                7 : begin
                    proc_path = "toe_top_toe_top.convert_axis_to_net_axis_512_3_U0";
                end
                8 : begin
                    proc_path = "toe_top_toe_top.convert_net_axis_to_axis_512_3_U0";
                end
                9 : begin
                    proc_path = "toe_top_toe_top.lookupReplyHandler_U0";
                end
                10 : begin
                    proc_path = "toe_top_toe_top.updateRequestSender_U0";
                end
                11 : begin
                    proc_path = "toe_top_toe_top.sessionIdManager_U0";
                end
                12 : begin
                    proc_path = "toe_top_toe_top.updateReplyHandler_U0";
                end
                13 : begin
                    proc_path = "toe_top_toe_top.reverseLookupTableInterface_U0";
                end
                14 : begin
                    proc_path = "toe_top_toe_top.state_table_U0";
                end
                15 : begin
                    proc_path = "toe_top_toe_top.rx_sar_table_U0";
                end
                16 : begin
                    proc_path = "toe_top_toe_top.tx_sar_table_U0";
                end
                17 : begin
                    proc_path = "toe_top_toe_top.listening_port_table_U0";
                end
                18 : begin
                    proc_path = "toe_top_toe_top.free_port_table_U0";
                end
                19 : begin
                    proc_path = "toe_top_toe_top.check_in_multiplexer_U0";
                end
                20 : begin
                    proc_path = "toe_top_toe_top.check_out_multiplexer_U0";
                end
                21 : begin
                    proc_path = "toe_top_toe_top.stream_merger_event_U0";
                end
                22 : begin
                    proc_path = "toe_top_toe_top.retransmit_timer_U0";
                end
                23 : begin
                    proc_path = "toe_top_toe_top.probe_timer_U0";
                end
                24 : begin
                    proc_path = "toe_top_toe_top.close_timer_U0";
                end
                25 : begin
                    proc_path = "toe_top_toe_top.stream_merger_ap_uint_16_U0";
                end
                26 : begin
                    proc_path = "toe_top_toe_top.event_engine_U0";
                end
                27 : begin
                    proc_path = "toe_top_toe_top.ack_delay_U0";
                end
                28 : begin
                    proc_path = "toe_top_toe_top.toe_process_ipv4_512_U0";
                end
                29 : begin
                    proc_path = "toe_top_toe_top.drop_optional_ip_header_512_U0";
                end
                30 : begin
                    proc_path = "toe_top_toe_top.lshiftWordByOctet_512_2_U0";
                end
                31 : begin
                    proc_path = "toe_top_toe_top.constructPseudoHeader_512_U0";
                end
                32 : begin
                    proc_path = "toe_top_toe_top.prependPseudoHeader_512_U0";
                end
                33 : begin
                    proc_path = "toe_top_toe_top.two_complement_subchecksums_512_11_U0";
                end
                34 : begin
                    proc_path = "toe_top_toe_top.toe_check_ipv4_checksum_32_U0";
                end
                35 : begin
                    proc_path = "toe_top_toe_top.processPseudoHeader_512_U0";
                end
                36 : begin
                    proc_path = "toe_top_toe_top.rshiftWordByOctet_net_axis_512_512_3_U0";
                end
                37 : begin
                    proc_path = "toe_top_toe_top.drop_optional_header_fields_512_U0";
                end
                38 : begin
                    proc_path = "toe_top_toe_top.parse_optional_header_fields_U0";
                end
                39 : begin
                    proc_path = "toe_top_toe_top.merge_header_meta_U0";
                end
                40 : begin
                    proc_path = "toe_top_toe_top.rxMetadataHandler_U0";
                end
                41 : begin
                    proc_path = "toe_top_toe_top.rxTcpFSM_U0";
                end
                42 : begin
                    proc_path = "toe_top_toe_top.rxPackageDropper_512_U0";
                end
                43 : begin
                    proc_path = "toe_top_toe_top.rxEventMerger_U0";
                end
                44 : begin
                    proc_path = "toe_top_toe_top.metaLoader_U0";
                end
                45 : begin
                    proc_path = "toe_top_toe_top.txEngMemAccessBreakdown_U0";
                end
                46 : begin
                    proc_path = "toe_top_toe_top.tupleSplitter_U0";
                end
                47 : begin
                    proc_path = "toe_top_toe_top.read_data_stitching_512_U0";
                end
                48 : begin
                    proc_path = "toe_top_toe_top.read_data_arbiter_512_U0";
                end
                49 : begin
                    proc_path = "toe_top_toe_top.lshiftWordByOctet_512_51_U0";
                end
                50 : begin
                    proc_path = "toe_top_toe_top.pseudoHeaderConstructionNew_512_U0";
                end
                51 : begin
                    proc_path = "toe_top_toe_top.two_complement_subchecksums_512_22_U0";
                end
                52 : begin
                    proc_path = "toe_top_toe_top.finalize_ipv4_checksum_32_U0";
                end
                53 : begin
                    proc_path = "toe_top_toe_top.remove_pseudo_header_512_U0";
                end
                54 : begin
                    proc_path = "toe_top_toe_top.rshiftWordByOctet_net_axis_512_512_53_U0";
                end
                55 : begin
                    proc_path = "toe_top_toe_top.insert_checksum_512_U0";
                end
                56 : begin
                    proc_path = "toe_top_toe_top.lshiftWordByOctet_512_52_U0";
                end
                57 : begin
                    proc_path = "toe_top_toe_top.generate_ipv4_512_U0";
                end
                58 : begin
                    proc_path = "toe_top_toe_top.rx_app_stream_if_U0";
                end
                59 : begin
                    proc_path = "toe_top_toe_top.rxAppMemDataRead_512_U0";
                end
                60 : begin
                    proc_path = "toe_top_toe_top.rx_app_if_U0";
                end
                61 : begin
                    proc_path = "toe_top_toe_top.stream_merger_appNotification_U0";
                end
                62 : begin
                    proc_path = "toe_top_toe_top.txEventMerger_U0";
                end
                63 : begin
                    proc_path = "toe_top_toe_top.txAppStatusHandler_U0";
                end
                64 : begin
                    proc_path = "toe_top_toe_top.tasi_metaLoader_U0";
                end
                65 : begin
                    proc_path = "toe_top_toe_top.toe_duplicate_stream_net_axis_512_U0";
                end
                66 : begin
                    proc_path = "toe_top_toe_top.tasi_pkg_pusher_512_U0";
                end
                67 : begin
                    proc_path = "toe_top_toe_top.tx_app_if_U0";
                end
                68 : begin
                    proc_path = "toe_top_toe_top.tx_app_table_U0";
                end
                default : begin
                    proc_path = "unknown";
                end
            endcase
        end
    endfunction

    // print the headlines of deadlock detection
    task print_dl_head;
        begin
            $display("\n//////////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", $time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            fp = $fopen("deadlock_db.dat", "w");
        end
    endtask

    // print the start of a cycle
    task print_cycle_start(input reg [488:0] proc_path, input integer cycle_id);
        begin
            $display("/////////////////////////");
            $display("// Dependence cycle %0d:", cycle_id);
            $display("// (1): Process: %0s", proc_path);
            $fdisplay(fp, "Dependence_Cycle_ID %0d", cycle_id);
            $fdisplay(fp, "Dependence_Process_ID 1");
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print the end of deadlock detection
    task print_dl_end(input integer num, input integer record_time);
        begin
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// Totally %0d cycles detected!", num);
            $display("////////////////////////////////////////////////////////////////////////");
            $display("// ERROR!!! DEADLOCK DETECTED at %0t ns! SIMULATION WILL BE STOPPED! //", record_time);
            $display("//////////////////////////////////////////////////////////////////////////////");
            $fdisplay(fp, "Dependence_Cycle_Number %0d", num);
            $fclose(fp);
        end
    endtask

    // print one proc component in the cycle
    task print_cycle_proc_comp(input reg [488:0] proc_path, input integer cycle_comp_id);
        begin
            $display("// (%0d): Process: %0s", cycle_comp_id, proc_path);
            $fdisplay(fp, "Dependence_Process_ID %0d", cycle_comp_id);
            $fdisplay(fp, "Dependence_Process_path %0s", proc_path);
        end
    endtask

    // print one channel component in the cycle
    task print_cycle_chan_comp(input [PROC_NUM - 1:0] dl_vec1, input [PROC_NUM - 1:0] dl_vec2);
        reg [456:0] chan_path;
        integer index1;
        integer index2;
        begin
            index1 = proc_index(dl_vec1);
            index2 = proc_index(dl_vec2);
            case (index1)
                0 : begin
                    case(index2)
                    41: begin
                        if (~entry_proc_U0.axis_data_count_c_blk_n) begin
                            if (~axis_data_count_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.axis_data_count_c_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.axis_data_count_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~axis_data_count_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.axis_data_count_c_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.axis_data_count_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~entry_proc_U0.axis_max_data_count_c_blk_n) begin
                            if (~axis_max_data_count_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.axis_max_data_count_c_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.axis_max_data_count_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~axis_max_data_count_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.axis_max_data_count_c_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.axis_max_data_count_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~entry_proc_U0.myIpAddress_c143_blk_n) begin
                            if (~myIpAddress_c143_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.myIpAddress_c143_U' written by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.myIpAddress_c143_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~myIpAddress_c143_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.myIpAddress_c143_U' read by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.myIpAddress_c143_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                1 : begin
                    case(index2)
                    28: begin
                        if (~convert_axis_to_net_axis_512_U0.ipRxData_internal_blk_n) begin
                            if (~ipRxData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.ipRxData_internal_U' written by process 'toe_top_toe_top.toe_process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ipRxData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~ipRxData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.ipRxData_internal_U' read by process 'toe_top_toe_top.toe_process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ipRxData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                2 : begin
                    case(index2)
                    59: begin
                        if (~convert_axis_to_net_axis_512_1_U0.rxBufferReadData_internal_blk_n) begin
                            if (~rxBufferReadData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxBufferReadData_internal_U' written by process 'toe_top_toe_top.rxAppMemDataRead_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferReadData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxBufferReadData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxBufferReadData_internal_U' read by process 'toe_top_toe_top.rxAppMemDataRead_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferReadData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                3 : begin
                    case(index2)
                    47: begin
                        if (~convert_axis_to_net_axis_512_2_U0.txBufferReadData_internal_blk_n) begin
                            if (~txBufferReadData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txBufferReadData_internal_U' written by process 'toe_top_toe_top.read_data_stitching_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferReadData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txBufferReadData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txBufferReadData_internal_U' read by process 'toe_top_toe_top.read_data_stitching_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferReadData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                4 : begin
                    case(index2)
                    57: begin
                        if (~convert_net_axis_to_axis_512_U0.ipTxData_internal_blk_n) begin
                            if (~ipTxData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.ipTxData_internal_U' written by process 'toe_top_toe_top.generate_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ipTxData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~ipTxData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.ipTxData_internal_U' read by process 'toe_top_toe_top.generate_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ipTxData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                5 : begin
                    case(index2)
                    42: begin
                        if (~convert_net_axis_to_axis_512_1_U0.rxBufferWriteData_internal_blk_n) begin
                            if (~rxBufferWriteData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxBufferWriteData_internal_U' written by process 'toe_top_toe_top.rxPackageDropper_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferWriteData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxBufferWriteData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxBufferWriteData_internal_U' read by process 'toe_top_toe_top.rxPackageDropper_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferWriteData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                6 : begin
                    case(index2)
                    66: begin
                        if (~convert_net_axis_to_axis_512_2_U0.txBufferWriteData_internal_blk_n) begin
                            if (~txBufferWriteData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txBufferWriteData_internal_U' written by process 'toe_top_toe_top.tasi_pkg_pusher_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferWriteData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txBufferWriteData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txBufferWriteData_internal_U' read by process 'toe_top_toe_top.tasi_pkg_pusher_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferWriteData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                7 : begin
                    case(index2)
                    65: begin
                        if (~convert_axis_to_net_axis_512_3_U0.txDataReq_internal_blk_n) begin
                            if (~txDataReq_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txDataReq_internal_U' written by process 'toe_top_toe_top.toe_duplicate_stream_net_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txDataReq_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txDataReq_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txDataReq_internal_U' read by process 'toe_top_toe_top.toe_duplicate_stream_net_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txDataReq_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                8 : begin
                    case(index2)
                    59: begin
                        if (~convert_net_axis_to_axis_512_3_U0.rxDataRsp_internal_blk_n) begin
                            if (~rxDataRsp_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxDataRsp_internal_U' written by process 'toe_top_toe_top.rxAppMemDataRead_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxDataRsp_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxDataRsp_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxDataRsp_internal_U' read by process 'toe_top_toe_top.rxAppMemDataRead_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxDataRsp_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                9 : begin
                    case(index2)
                    67: begin
                        if (~lookupReplyHandler_U0.txApp2sLookup_req_blk_n) begin
                            if (~txApp2sLookup_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2sLookup_req_U' written by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2sLookup_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2sLookup_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2sLookup_req_U' read by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2sLookup_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~lookupReplyHandler_U0.sLookup2txApp_rsp_blk_n) begin
                            if (~sLookup2txApp_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sLookup2txApp_rsp_U' written by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2txApp_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sLookup2txApp_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sLookup2txApp_rsp_U' read by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2txApp_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    40: begin
                        if (~lookupReplyHandler_U0.rxEng2sLookup_req_blk_n) begin
                            if (~rxEng2sLookup_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2sLookup_req_U' written by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2sLookup_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2sLookup_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2sLookup_req_U' read by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2sLookup_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~lookupReplyHandler_U0.sLookup2rxEng_rsp_blk_n) begin
                            if (~sLookup2rxEng_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sLookup2rxEng_rsp_U' written by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2rxEng_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sLookup2rxEng_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sLookup2rxEng_rsp_U' read by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2rxEng_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    11: begin
                        if (~lookupReplyHandler_U0.slc_sessionIdFreeList_blk_n) begin
                            if (~slc_sessionIdFreeList_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.slc_sessionIdFreeList_U' written by process 'toe_top_toe_top.sessionIdManager_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionIdFreeList_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~slc_sessionIdFreeList_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.slc_sessionIdFreeList_U' read by process 'toe_top_toe_top.sessionIdManager_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionIdFreeList_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    10: begin
                        if (~lookupReplyHandler_U0.sessionInsert_req_blk_n) begin
                            if (~sessionInsert_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sessionInsert_req_U' written by process 'toe_top_toe_top.updateRequestSender_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sessionInsert_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sessionInsert_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sessionInsert_req_U' read by process 'toe_top_toe_top.updateRequestSender_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sessionInsert_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    12: begin
                        if (~lookupReplyHandler_U0.slc_sessionInsert_rsp_blk_n) begin
                            if (~slc_sessionInsert_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.slc_sessionInsert_rsp_U' written by process 'toe_top_toe_top.updateReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionInsert_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~slc_sessionInsert_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.slc_sessionInsert_rsp_U' read by process 'toe_top_toe_top.updateReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionInsert_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~lookupReplyHandler_U0.reverseLupInsertFifo_blk_n) begin
                            if (~reverseLupInsertFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.reverseLupInsertFifo_U' written by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.reverseLupInsertFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~reverseLupInsertFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.reverseLupInsertFifo_U' read by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.reverseLupInsertFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                10 : begin
                    case(index2)
                    9: begin
                        if (~updateRequestSender_U0.sessionInsert_req_blk_n) begin
                            if (~sessionInsert_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sessionInsert_req_U' written by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sessionInsert_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sessionInsert_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sessionInsert_req_U' read by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sessionInsert_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~updateRequestSender_U0.sessionDelete_req_blk_n) begin
                            if (~sessionDelete_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sessionDelete_req_U' written by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sessionDelete_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sessionDelete_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sessionDelete_req_U' read by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sessionDelete_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    11: begin
                        if (~updateRequestSender_U0.slc_sessionIdFinFifo_blk_n) begin
                            if (~slc_sessionIdFinFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.slc_sessionIdFinFifo_U' written by process 'toe_top_toe_top.sessionIdManager_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionIdFinFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~slc_sessionIdFinFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.slc_sessionIdFinFifo_U' read by process 'toe_top_toe_top.sessionIdManager_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionIdFinFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                11 : begin
                    case(index2)
                    10: begin
                        if (~sessionIdManager_U0.slc_sessionIdFinFifo_blk_n) begin
                            if (~slc_sessionIdFinFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.slc_sessionIdFinFifo_U' written by process 'toe_top_toe_top.updateRequestSender_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionIdFinFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~slc_sessionIdFinFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.slc_sessionIdFinFifo_U' read by process 'toe_top_toe_top.updateRequestSender_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionIdFinFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    9: begin
                        if (~sessionIdManager_U0.slc_sessionIdFreeList_blk_n) begin
                            if (~slc_sessionIdFreeList_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.slc_sessionIdFreeList_U' written by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionIdFreeList_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~slc_sessionIdFreeList_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.slc_sessionIdFreeList_U' read by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionIdFreeList_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                12 : begin
                    case(index2)
                    9: begin
                        if (~updateReplyHandler_U0.slc_sessionInsert_rsp_blk_n) begin
                            if (~slc_sessionInsert_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.slc_sessionInsert_rsp_U' written by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionInsert_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~slc_sessionInsert_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.slc_sessionInsert_rsp_U' read by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.slc_sessionInsert_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                13 : begin
                    case(index2)
                    0: begin
                        if (~reverseLookupTableInterface_U0.myIpAddress_blk_n) begin
                            if (~myIpAddress_c143_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.myIpAddress_c143_U' written by process 'toe_top_toe_top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.myIpAddress_c143_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~myIpAddress_c143_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.myIpAddress_c143_U' read by process 'toe_top_toe_top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.myIpAddress_c143_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    67: begin
                        if (~reverseLookupTableInterface_U0.myIpAddress_c_blk_n) begin
                            if (~myIpAddress_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.myIpAddress_c_U' written by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.myIpAddress_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~myIpAddress_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.myIpAddress_c_U' read by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.myIpAddress_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    9: begin
                        if (~reverseLookupTableInterface_U0.reverseLupInsertFifo_blk_n) begin
                            if (~reverseLupInsertFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.reverseLupInsertFifo_U' written by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.reverseLupInsertFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~reverseLupInsertFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.reverseLupInsertFifo_U' read by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.reverseLupInsertFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~reverseLookupTableInterface_U0.stateTable2sLookup_releaseSession_blk_n) begin
                            if (~stateTable2sLookup_releaseSession_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.stateTable2sLookup_releaseSession_U' written by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2sLookup_releaseSession_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2sLookup_releaseSession_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.stateTable2sLookup_releaseSession_U' read by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2sLookup_releaseSession_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    18: begin
                        if (~reverseLookupTableInterface_U0.sLookup2portTable_releasePort_blk_n) begin
                            if (~sLookup2portTable_releasePort_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sLookup2portTable_releasePort_U' written by process 'toe_top_toe_top.free_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2portTable_releasePort_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sLookup2portTable_releasePort_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sLookup2portTable_releasePort_U' read by process 'toe_top_toe_top.free_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2portTable_releasePort_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    10: begin
                        if (~reverseLookupTableInterface_U0.sessionDelete_req_blk_n) begin
                            if (~sessionDelete_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sessionDelete_req_U' written by process 'toe_top_toe_top.updateRequestSender_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sessionDelete_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sessionDelete_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sessionDelete_req_U' read by process 'toe_top_toe_top.updateRequestSender_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sessionDelete_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    44: begin
                        if (~reverseLookupTableInterface_U0.txEng2sLookup_rev_req_blk_n) begin
                            if (~txEng2sLookup_rev_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng2sLookup_rev_req_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2sLookup_rev_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng2sLookup_rev_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng2sLookup_rev_req_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2sLookup_rev_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    46: begin
                        if (~reverseLookupTableInterface_U0.sLookup2txEng_rev_rsp_blk_n) begin
                            if (~sLookup2txEng_rev_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sLookup2txEng_rev_rsp_U' written by process 'toe_top_toe_top.tupleSplitter_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2txEng_rev_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sLookup2txEng_rev_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sLookup2txEng_rev_rsp_U' read by process 'toe_top_toe_top.tupleSplitter_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2txEng_rev_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                14 : begin
                    case(index2)
                    67: begin
                        if (~state_table_U0.txApp2stateTable_upd_req_blk_n) begin
                            if (~txApp2stateTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2stateTable_upd_req_U' written by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2stateTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2stateTable_upd_req_U' read by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~state_table_U0.stateTable2txApp_upd_rsp_blk_n) begin
                            if (~stateTable2txApp_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.stateTable2txApp_upd_rsp_U' written by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2txApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2txApp_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.stateTable2txApp_upd_rsp_U' read by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2txApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    64: begin
                        if (~state_table_U0.txApp2stateTable_req_blk_n) begin
                            if (~txApp2stateTable_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2stateTable_req_U' written by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2stateTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2stateTable_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2stateTable_req_U' read by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2stateTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~state_table_U0.stateTable2txApp_rsp_blk_n) begin
                            if (~stateTable2txApp_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.stateTable2txApp_rsp_U' written by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2txApp_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2txApp_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.stateTable2txApp_rsp_U' read by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2txApp_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    41: begin
                        if (~state_table_U0.rxEng2stateTable_upd_req_blk_n) begin
                            if (~rxEng2stateTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2stateTable_upd_req_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2stateTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2stateTable_upd_req_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~state_table_U0.stateTable2rxEng_upd_rsp_blk_n) begin
                            if (~stateTable2rxEng_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.stateTable2rxEng_upd_rsp_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2rxEng_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.stateTable2rxEng_upd_rsp_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~state_table_U0.stateTable2sLookup_releaseSession_blk_n) begin
                            if (~stateTable2sLookup_releaseSession_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.stateTable2sLookup_releaseSession_U' written by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2sLookup_releaseSession_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2sLookup_releaseSession_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.stateTable2sLookup_releaseSession_U' read by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2sLookup_releaseSession_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    25: begin
                        if (~state_table_U0.timer2stateTable_releaseState_blk_n) begin
                            if (~timer2stateTable_releaseState_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.timer2stateTable_releaseState_U' written by process 'toe_top_toe_top.stream_merger_ap_uint_16_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~timer2stateTable_releaseState_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.timer2stateTable_releaseState_U' read by process 'toe_top_toe_top.stream_merger_ap_uint_16_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                15 : begin
                    case(index2)
                    44: begin
                        if (~rx_sar_table_U0.txEng2rxSar_req_blk_n) begin
                            if (~txEng2rxSar_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng2rxSar_req_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2rxSar_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng2rxSar_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng2rxSar_req_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2rxSar_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rx_sar_table_U0.rxSar2txEng_rsp_blk_n) begin
                            if (~rxSar2txEng_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxSar2txEng_rsp_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2txEng_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxSar2txEng_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxSar2txEng_rsp_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2txEng_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    58: begin
                        if (~rx_sar_table_U0.rxApp2rxSar_upd_req_blk_n) begin
                            if (~rxApp2rxSar_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxApp2rxSar_upd_req_U' written by process 'toe_top_toe_top.rx_app_stream_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxApp2rxSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxApp2rxSar_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxApp2rxSar_upd_req_U' read by process 'toe_top_toe_top.rx_app_stream_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxApp2rxSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rx_sar_table_U0.rxSar2rxApp_upd_rsp_blk_n) begin
                            if (~rxSar2rxApp_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxSar2rxApp_upd_rsp_U' written by process 'toe_top_toe_top.rx_app_stream_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2rxApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxSar2rxApp_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxSar2rxApp_upd_rsp_U' read by process 'toe_top_toe_top.rx_app_stream_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2rxApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    41: begin
                        if (~rx_sar_table_U0.rxEng2rxSar_upd_req_blk_n) begin
                            if (~rxEng2rxSar_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2rxSar_upd_req_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2rxSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2rxSar_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2rxSar_upd_req_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2rxSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rx_sar_table_U0.rxSar2rxEng_upd_rsp_blk_n) begin
                            if (~rxSar2rxEng_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxSar2rxEng_upd_rsp_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxSar2rxEng_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxSar2rxEng_upd_rsp_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                16 : begin
                    case(index2)
                    44: begin
                        if (~tx_sar_table_U0.txEng2txSar_upd_req_blk_n) begin
                            if (~txEng2txSar_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng2txSar_upd_req_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng2txSar_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng2txSar_upd_req_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~tx_sar_table_U0.txSar2txEng_upd_rsp_blk_n) begin
                            if (~txSar2txEng_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txSar2txEng_upd_rsp_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txSar2txEng_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txSar2txEng_upd_rsp_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    68: begin
                        if (~tx_sar_table_U0.txSar2txApp_ack_push_blk_n) begin
                            if (~txSar2txApp_ack_push_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txSar2txApp_ack_push_U' written by process 'toe_top_toe_top.tx_app_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txApp_ack_push_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txSar2txApp_ack_push_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txSar2txApp_ack_push_U' read by process 'toe_top_toe_top.tx_app_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txApp_ack_push_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    63: begin
                        if (~tx_sar_table_U0.txApp2txSar_push_blk_n) begin
                            if (~txApp2txSar_push_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2txSar_push_U' written by process 'toe_top_toe_top.txAppStatusHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txSar_push_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2txSar_push_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2txSar_push_U' read by process 'toe_top_toe_top.txAppStatusHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txSar_push_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    41: begin
                        if (~tx_sar_table_U0.rxEng2txSar_upd_req_blk_n) begin
                            if (~rxEng2txSar_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2txSar_upd_req_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2txSar_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2txSar_upd_req_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~tx_sar_table_U0.txSar2rxEng_upd_rsp_blk_n) begin
                            if (~txSar2rxEng_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txSar2rxEng_upd_rsp_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txSar2rxEng_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txSar2rxEng_upd_rsp_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                17 : begin
                    case(index2)
                    60: begin
                        if (~listening_port_table_U0.rxApp2portTable_listen_req_blk_n) begin
                            if (~rxApp2portTable_listen_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxApp2portTable_listen_req_U' written by process 'toe_top_toe_top.rx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxApp2portTable_listen_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxApp2portTable_listen_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxApp2portTable_listen_req_U' read by process 'toe_top_toe_top.rx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxApp2portTable_listen_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~listening_port_table_U0.portTable2rxApp_listen_rsp_blk_n) begin
                            if (~portTable2rxApp_listen_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.portTable2rxApp_listen_rsp_U' written by process 'toe_top_toe_top.rx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2rxApp_listen_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~portTable2rxApp_listen_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.portTable2rxApp_listen_rsp_U' read by process 'toe_top_toe_top.rx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2rxApp_listen_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (~listening_port_table_U0.pt_portCheckListening_req_fifo_blk_n) begin
                            if (~pt_portCheckListening_req_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.pt_portCheckListening_req_fifo_U' written by process 'toe_top_toe_top.check_in_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckListening_req_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~pt_portCheckListening_req_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.pt_portCheckListening_req_fifo_U' read by process 'toe_top_toe_top.check_in_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckListening_req_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (~listening_port_table_U0.pt_portCheckListening_rsp_fifo_blk_n) begin
                            if (~pt_portCheckListening_rsp_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.pt_portCheckListening_rsp_fifo_U' written by process 'toe_top_toe_top.check_out_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckListening_rsp_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~pt_portCheckListening_rsp_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.pt_portCheckListening_rsp_fifo_U' read by process 'toe_top_toe_top.check_out_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckListening_rsp_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                18 : begin
                    case(index2)
                    13: begin
                        if (~free_port_table_U0.sLookup2portTable_releasePort_blk_n) begin
                            if (~sLookup2portTable_releasePort_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sLookup2portTable_releasePort_U' written by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2portTable_releasePort_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sLookup2portTable_releasePort_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sLookup2portTable_releasePort_U' read by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2portTable_releasePort_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (~free_port_table_U0.pt_portCheckUsed_req_fifo_blk_n) begin
                            if (~pt_portCheckUsed_req_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.pt_portCheckUsed_req_fifo_U' written by process 'toe_top_toe_top.check_in_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckUsed_req_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~pt_portCheckUsed_req_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.pt_portCheckUsed_req_fifo_U' read by process 'toe_top_toe_top.check_in_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckUsed_req_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (~free_port_table_U0.pt_portCheckUsed_rsp_fifo_blk_n) begin
                            if (~pt_portCheckUsed_rsp_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.pt_portCheckUsed_rsp_fifo_U' written by process 'toe_top_toe_top.check_out_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckUsed_rsp_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~pt_portCheckUsed_rsp_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.pt_portCheckUsed_rsp_fifo_U' read by process 'toe_top_toe_top.check_out_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckUsed_rsp_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    67: begin
                        if (~free_port_table_U0.portTable2txApp_port_rsp_blk_n) begin
                            if (~portTable2txApp_port_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.portTable2txApp_port_rsp_U' written by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2txApp_port_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~portTable2txApp_port_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.portTable2txApp_port_rsp_U' read by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2txApp_port_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                19 : begin
                    case(index2)
                    35: begin
                        if (~check_in_multiplexer_U0.rxEng2portTable_check_req_blk_n) begin
                            if (~rxEng2portTable_check_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2portTable_check_req_U' written by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2portTable_check_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2portTable_check_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2portTable_check_req_U' read by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2portTable_check_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    17: begin
                        if (~check_in_multiplexer_U0.pt_portCheckListening_req_fifo_blk_n) begin
                            if (~pt_portCheckListening_req_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.pt_portCheckListening_req_fifo_U' written by process 'toe_top_toe_top.listening_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckListening_req_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~pt_portCheckListening_req_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.pt_portCheckListening_req_fifo_U' read by process 'toe_top_toe_top.listening_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckListening_req_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (~check_in_multiplexer_U0.pt_dstFifo_blk_n) begin
                            if (~pt_dstFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.pt_dstFifo_U' written by process 'toe_top_toe_top.check_out_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_dstFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~pt_dstFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.pt_dstFifo_U' read by process 'toe_top_toe_top.check_out_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_dstFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    18: begin
                        if (~check_in_multiplexer_U0.pt_portCheckUsed_req_fifo_blk_n) begin
                            if (~pt_portCheckUsed_req_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.pt_portCheckUsed_req_fifo_U' written by process 'toe_top_toe_top.free_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckUsed_req_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~pt_portCheckUsed_req_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.pt_portCheckUsed_req_fifo_U' read by process 'toe_top_toe_top.free_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckUsed_req_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                20 : begin
                    case(index2)
                    19: begin
                        if (~check_out_multiplexer_U0.pt_dstFifo_blk_n) begin
                            if (~pt_dstFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.pt_dstFifo_U' written by process 'toe_top_toe_top.check_in_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_dstFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~pt_dstFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.pt_dstFifo_U' read by process 'toe_top_toe_top.check_in_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_dstFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    17: begin
                        if (~check_out_multiplexer_U0.pt_portCheckListening_rsp_fifo_blk_n) begin
                            if (~pt_portCheckListening_rsp_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.pt_portCheckListening_rsp_fifo_U' written by process 'toe_top_toe_top.listening_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckListening_rsp_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~pt_portCheckListening_rsp_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.pt_portCheckListening_rsp_fifo_U' read by process 'toe_top_toe_top.listening_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckListening_rsp_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    40: begin
                        if (~check_out_multiplexer_U0.portTable2rxEng_check_rsp_blk_n) begin
                            if (~portTable2rxEng_check_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.portTable2rxEng_check_rsp_U' written by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2rxEng_check_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~portTable2rxEng_check_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.portTable2rxEng_check_rsp_U' read by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2rxEng_check_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    18: begin
                        if (~check_out_multiplexer_U0.pt_portCheckUsed_rsp_fifo_blk_n) begin
                            if (~pt_portCheckUsed_rsp_fifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.pt_portCheckUsed_rsp_fifo_U' written by process 'toe_top_toe_top.free_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckUsed_rsp_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~pt_portCheckUsed_rsp_fifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.pt_portCheckUsed_rsp_fifo_U' read by process 'toe_top_toe_top.free_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.pt_portCheckUsed_rsp_fifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                21 : begin
                    case(index2)
                    22: begin
                        if (~stream_merger_event_U0.rtTimer2eventEng_setEvent_blk_n) begin
                            if (~rtTimer2eventEng_setEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rtTimer2eventEng_setEvent_U' written by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rtTimer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rtTimer2eventEng_setEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rtTimer2eventEng_setEvent_U' read by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rtTimer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    26: begin
                        if (~stream_merger_event_U0.timer2eventEng_setEvent_blk_n) begin
                            if (~timer2eventEng_setEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.timer2eventEng_setEvent_U' written by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~timer2eventEng_setEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.timer2eventEng_setEvent_U' read by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    23: begin
                        if (~stream_merger_event_U0.probeTimer2eventEng_setEvent_blk_n) begin
                            if (~probeTimer2eventEng_setEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.probeTimer2eventEng_setEvent_U' written by process 'toe_top_toe_top.probe_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.probeTimer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~probeTimer2eventEng_setEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.probeTimer2eventEng_setEvent_U' read by process 'toe_top_toe_top.probe_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.probeTimer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                22 : begin
                    case(index2)
                    41: begin
                        if (~retransmit_timer_U0.rxEng2timer_clearRetransmitTimer_blk_n) begin
                            if (~rxEng2timer_clearRetransmitTimer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2timer_clearRetransmitTimer_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_clearRetransmitTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2timer_clearRetransmitTimer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2timer_clearRetransmitTimer_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_clearRetransmitTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    44: begin
                        if (~retransmit_timer_U0.txEng2timer_setRetransmitTimer_blk_n) begin
                            if (~txEng2timer_setRetransmitTimer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng2timer_setRetransmitTimer_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2timer_setRetransmitTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng2timer_setRetransmitTimer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng2timer_setRetransmitTimer_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2timer_setRetransmitTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    21: begin
                        if (~retransmit_timer_U0.rtTimer2eventEng_setEvent_blk_n) begin
                            if (~rtTimer2eventEng_setEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rtTimer2eventEng_setEvent_U' written by process 'toe_top_toe_top.stream_merger_event_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rtTimer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rtTimer2eventEng_setEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rtTimer2eventEng_setEvent_U' read by process 'toe_top_toe_top.stream_merger_event_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rtTimer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    25: begin
                        if (~retransmit_timer_U0.rtTimer2stateTable_releaseState_blk_n) begin
                            if (~rtTimer2stateTable_releaseState_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rtTimer2stateTable_releaseState_U' written by process 'toe_top_toe_top.stream_merger_ap_uint_16_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rtTimer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rtTimer2stateTable_releaseState_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rtTimer2stateTable_releaseState_U' read by process 'toe_top_toe_top.stream_merger_ap_uint_16_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rtTimer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    67: begin
                        if (~retransmit_timer_U0.timer2txApp_notification_blk_n) begin
                            if (~timer2txApp_notification_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.timer2txApp_notification_U' written by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2txApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~timer2txApp_notification_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.timer2txApp_notification_U' read by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2txApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    61: begin
                        if (~retransmit_timer_U0.timer2rxApp_notification_blk_n) begin
                            if (~timer2rxApp_notification_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.timer2rxApp_notification_U' written by process 'toe_top_toe_top.stream_merger_appNotification_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2rxApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~timer2rxApp_notification_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.timer2rxApp_notification_U' read by process 'toe_top_toe_top.stream_merger_appNotification_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2rxApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                23 : begin
                    case(index2)
                    44: begin
                        if (~probe_timer_U0.txEng2timer_setProbeTimer_blk_n) begin
                            if (~txEng2timer_setProbeTimer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng2timer_setProbeTimer_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2timer_setProbeTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng2timer_setProbeTimer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng2timer_setProbeTimer_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2timer_setProbeTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    41: begin
                        if (~probe_timer_U0.rxEng2timer_clearProbeTimer_blk_n) begin
                            if (~rxEng2timer_clearProbeTimer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2timer_clearProbeTimer_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_clearProbeTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2timer_clearProbeTimer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2timer_clearProbeTimer_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_clearProbeTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    21: begin
                        if (~probe_timer_U0.probeTimer2eventEng_setEvent_blk_n) begin
                            if (~probeTimer2eventEng_setEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.probeTimer2eventEng_setEvent_U' written by process 'toe_top_toe_top.stream_merger_event_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.probeTimer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~probeTimer2eventEng_setEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.probeTimer2eventEng_setEvent_U' read by process 'toe_top_toe_top.stream_merger_event_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.probeTimer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                24 : begin
                    case(index2)
                    41: begin
                        if (~close_timer_U0.rxEng2timer_setCloseTimer_blk_n) begin
                            if (~rxEng2timer_setCloseTimer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2timer_setCloseTimer_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_setCloseTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2timer_setCloseTimer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2timer_setCloseTimer_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_setCloseTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    25: begin
                        if (~close_timer_U0.closeTimer2stateTable_releaseState_blk_n) begin
                            if (~closeTimer2stateTable_releaseState_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.closeTimer2stateTable_releaseState_U' written by process 'toe_top_toe_top.stream_merger_ap_uint_16_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.closeTimer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~closeTimer2stateTable_releaseState_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.closeTimer2stateTable_releaseState_U' read by process 'toe_top_toe_top.stream_merger_ap_uint_16_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.closeTimer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                25 : begin
                    case(index2)
                    24: begin
                        if (~stream_merger_ap_uint_16_U0.closeTimer2stateTable_releaseState_blk_n) begin
                            if (~closeTimer2stateTable_releaseState_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.closeTimer2stateTable_releaseState_U' written by process 'toe_top_toe_top.close_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.closeTimer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~closeTimer2stateTable_releaseState_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.closeTimer2stateTable_releaseState_U' read by process 'toe_top_toe_top.close_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.closeTimer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~stream_merger_ap_uint_16_U0.timer2stateTable_releaseState_blk_n) begin
                            if (~timer2stateTable_releaseState_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.timer2stateTable_releaseState_U' written by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~timer2stateTable_releaseState_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.timer2stateTable_releaseState_U' read by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    22: begin
                        if (~stream_merger_ap_uint_16_U0.rtTimer2stateTable_releaseState_blk_n) begin
                            if (~rtTimer2stateTable_releaseState_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rtTimer2stateTable_releaseState_U' written by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rtTimer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rtTimer2stateTable_releaseState_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rtTimer2stateTable_releaseState_U' read by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rtTimer2stateTable_releaseState_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                26 : begin
                    case(index2)
                    43: begin
                        if (~event_engine_U0.rxEng2eventEng_setEvent_blk_n) begin
                            if (~rxEng2eventEng_setEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2eventEng_setEvent_U' written by process 'toe_top_toe_top.rxEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2eventEng_setEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2eventEng_setEvent_U' read by process 'toe_top_toe_top.rxEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    27: begin
                        if (~event_engine_U0.eventEng2ackDelay_event_blk_n) begin
                            if (~eventEng2ackDelay_event_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.eventEng2ackDelay_event_U' written by process 'toe_top_toe_top.ack_delay_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.eventEng2ackDelay_event_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~eventEng2ackDelay_event_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.eventEng2ackDelay_event_U' read by process 'toe_top_toe_top.ack_delay_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.eventEng2ackDelay_event_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~event_engine_U0.ackDelayFifoReadCount_blk_n) begin
                            if (~ackDelayFifoReadCount_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.ackDelayFifoReadCount_U' written by process 'toe_top_toe_top.ack_delay_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ackDelayFifoReadCount_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~ackDelayFifoReadCount_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.ackDelayFifoReadCount_U' read by process 'toe_top_toe_top.ack_delay_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ackDelayFifoReadCount_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~event_engine_U0.ackDelayFifoWriteCount_blk_n) begin
                            if (~ackDelayFifoWriteCount_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.ackDelayFifoWriteCount_U' written by process 'toe_top_toe_top.ack_delay_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ackDelayFifoWriteCount_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~ackDelayFifoWriteCount_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.ackDelayFifoWriteCount_U' read by process 'toe_top_toe_top.ack_delay_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ackDelayFifoWriteCount_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    21: begin
                        if (~event_engine_U0.timer2eventEng_setEvent_blk_n) begin
                            if (~timer2eventEng_setEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.timer2eventEng_setEvent_U' written by process 'toe_top_toe_top.stream_merger_event_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~timer2eventEng_setEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.timer2eventEng_setEvent_U' read by process 'toe_top_toe_top.stream_merger_event_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    62: begin
                        if (~event_engine_U0.txApp2eventEng_setEvent_blk_n) begin
                            if (~txApp2eventEng_setEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2eventEng_setEvent_U' written by process 'toe_top_toe_top.txEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2eventEng_setEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2eventEng_setEvent_U' read by process 'toe_top_toe_top.txEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    44: begin
                        if (~event_engine_U0.txEngFifoReadCount_blk_n) begin
                            if (~txEngFifoReadCount_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEngFifoReadCount_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEngFifoReadCount_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEngFifoReadCount_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEngFifoReadCount_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEngFifoReadCount_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                27 : begin
                    case(index2)
                    26: begin
                        if (~ack_delay_U0.eventEng2ackDelay_event_blk_n) begin
                            if (~eventEng2ackDelay_event_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.eventEng2ackDelay_event_U' written by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.eventEng2ackDelay_event_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~eventEng2ackDelay_event_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.eventEng2ackDelay_event_U' read by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.eventEng2ackDelay_event_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~ack_delay_U0.ackDelayFifoReadCount_blk_n) begin
                            if (~ackDelayFifoReadCount_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.ackDelayFifoReadCount_U' written by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ackDelayFifoReadCount_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~ackDelayFifoReadCount_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.ackDelayFifoReadCount_U' read by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ackDelayFifoReadCount_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~ack_delay_U0.ackDelayFifoWriteCount_blk_n) begin
                            if (~ackDelayFifoWriteCount_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.ackDelayFifoWriteCount_U' written by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ackDelayFifoWriteCount_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~ackDelayFifoWriteCount_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.ackDelayFifoWriteCount_U' read by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ackDelayFifoWriteCount_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    44: begin
                        if (~ack_delay_U0.eventEng2txEng_event_blk_n) begin
                            if (~eventEng2txEng_event_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.eventEng2txEng_event_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.eventEng2txEng_event_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~eventEng2txEng_event_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.eventEng2txEng_event_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.eventEng2txEng_event_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                28 : begin
                    case(index2)
                    1: begin
                        if (~toe_process_ipv4_512_U0.ipRxData_internal_blk_n) begin
                            if (~ipRxData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.ipRxData_internal_U' written by process 'toe_top_toe_top.convert_axis_to_net_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ipRxData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~ipRxData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.ipRxData_internal_U' read by process 'toe_top_toe_top.convert_axis_to_net_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ipRxData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    29: begin
                        if (~toe_process_ipv4_512_U0.rxEng_dataBuffer0_blk_n) begin
                            if (~rxEng_dataBuffer0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer0_U' written by process 'toe_top_toe_top.drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer0_U' read by process 'toe_top_toe_top.drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~toe_process_ipv4_512_U0.rx_process2dropLengthFifo_blk_n) begin
                            if (~rx_process2dropLengthFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rx_process2dropLengthFifo_U' written by process 'toe_top_toe_top.drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rx_process2dropLengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_process2dropLengthFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rx_process2dropLengthFifo_U' read by process 'toe_top_toe_top.drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rx_process2dropLengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    31: begin
                        if (~toe_process_ipv4_512_U0.rxEng_ipMetaFifo_blk_n) begin
                            if (~rxEng_ipMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_ipMetaFifo_U' written by process 'toe_top_toe_top.constructPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_ipMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_ipMetaFifo_U' read by process 'toe_top_toe_top.constructPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                29 : begin
                    case(index2)
                    28: begin
                        if (~drop_optional_ip_header_512_U0.rx_process2dropLengthFifo_blk_n) begin
                            if (~rx_process2dropLengthFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rx_process2dropLengthFifo_U' written by process 'toe_top_toe_top.toe_process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rx_process2dropLengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rx_process2dropLengthFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rx_process2dropLengthFifo_U' read by process 'toe_top_toe_top.toe_process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rx_process2dropLengthFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~drop_optional_ip_header_512_U0.rxEng_dataBuffer0_blk_n) begin
                            if (~rxEng_dataBuffer0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer0_U' written by process 'toe_top_toe_top.toe_process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer0_U' read by process 'toe_top_toe_top.toe_process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    30: begin
                        if (~drop_optional_ip_header_512_U0.rxEng_dataBuffer4_blk_n) begin
                            if (~rxEng_dataBuffer4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer4_U' written by process 'toe_top_toe_top.lshiftWordByOctet_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer4_U' read by process 'toe_top_toe_top.lshiftWordByOctet_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                30 : begin
                    case(index2)
                    32: begin
                        if (~lshiftWordByOctet_512_2_U0.rxEng_dataBuffer5_blk_n) begin
                            if (~rxEng_dataBuffer5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer5_U' written by process 'toe_top_toe_top.prependPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer5_U' read by process 'toe_top_toe_top.prependPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    29: begin
                        if (~lshiftWordByOctet_512_2_U0.rxEng_dataBuffer4_blk_n) begin
                            if (~rxEng_dataBuffer4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer4_U' written by process 'toe_top_toe_top.drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer4_U' read by process 'toe_top_toe_top.drop_optional_ip_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                31 : begin
                    case(index2)
                    28: begin
                        if (~constructPseudoHeader_512_U0.rxEng_ipMetaFifo_blk_n) begin
                            if (~rxEng_ipMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_ipMetaFifo_U' written by process 'toe_top_toe_top.toe_process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_ipMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_ipMetaFifo_U' read by process 'toe_top_toe_top.toe_process_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    32: begin
                        if (~constructPseudoHeader_512_U0.rxEng_pseudoHeaderFifo_blk_n) begin
                            if (~rxEng_pseudoHeaderFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_pseudoHeaderFifo_U' written by process 'toe_top_toe_top.prependPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_pseudoHeaderFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_pseudoHeaderFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_pseudoHeaderFifo_U' read by process 'toe_top_toe_top.prependPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_pseudoHeaderFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                32 : begin
                    case(index2)
                    31: begin
                        if (~prependPseudoHeader_512_U0.rxEng_pseudoHeaderFifo_blk_n) begin
                            if (~rxEng_pseudoHeaderFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_pseudoHeaderFifo_U' written by process 'toe_top_toe_top.constructPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_pseudoHeaderFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_pseudoHeaderFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_pseudoHeaderFifo_U' read by process 'toe_top_toe_top.constructPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_pseudoHeaderFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    33: begin
                        if (~prependPseudoHeader_512_U0.rxEng_dataBuffer1_blk_n) begin
                            if (~rxEng_dataBuffer1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer1_U' written by process 'toe_top_toe_top.two_complement_subchecksums_512_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer1_U' read by process 'toe_top_toe_top.two_complement_subchecksums_512_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    30: begin
                        if (~prependPseudoHeader_512_U0.rxEng_dataBuffer5_blk_n) begin
                            if (~rxEng_dataBuffer5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer5_U' written by process 'toe_top_toe_top.lshiftWordByOctet_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer5_U' read by process 'toe_top_toe_top.lshiftWordByOctet_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                33 : begin
                    case(index2)
                    32: begin
                        if (~two_complement_subchecksums_512_11_U0.rxEng_dataBuffer1_blk_n) begin
                            if (~rxEng_dataBuffer1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer1_U' written by process 'toe_top_toe_top.prependPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer1_U' read by process 'toe_top_toe_top.prependPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    35: begin
                        if (~two_complement_subchecksums_512_11_U0.rxEng_dataBuffer2_blk_n) begin
                            if (~rxEng_dataBuffer2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer2_U' written by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer2_U' read by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    34: begin
                        if (~two_complement_subchecksums_512_11_U0.subSumFifo_blk_n) begin
                            if (~subSumFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.subSumFifo_U' written by process 'toe_top_toe_top.toe_check_ipv4_checksum_32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.subSumFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~subSumFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.subSumFifo_U' read by process 'toe_top_toe_top.toe_check_ipv4_checksum_32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.subSumFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                34 : begin
                    case(index2)
                    33: begin
                        if (~toe_check_ipv4_checksum_32_U0.subSumFifo_blk_n) begin
                            if (~subSumFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.subSumFifo_U' written by process 'toe_top_toe_top.two_complement_subchecksums_512_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.subSumFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~subSumFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.subSumFifo_U' read by process 'toe_top_toe_top.two_complement_subchecksums_512_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.subSumFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    35: begin
                        if (~toe_check_ipv4_checksum_32_U0.rxEng_checksumValidFifo_blk_n) begin
                            if (~rxEng_checksumValidFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_checksumValidFifo_U' written by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_checksumValidFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_checksumValidFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_checksumValidFifo_U' read by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_checksumValidFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                35 : begin
                    case(index2)
                    33: begin
                        if (~processPseudoHeader_512_U0.rxEng_dataBuffer2_blk_n) begin
                            if (~rxEng_dataBuffer2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer2_U' written by process 'toe_top_toe_top.two_complement_subchecksums_512_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer2_U' read by process 'toe_top_toe_top.two_complement_subchecksums_512_11_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    34: begin
                        if (~processPseudoHeader_512_U0.rxEng_checksumValidFifo_blk_n) begin
                            if (~rxEng_checksumValidFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_checksumValidFifo_U' written by process 'toe_top_toe_top.toe_check_ipv4_checksum_32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_checksumValidFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_checksumValidFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_checksumValidFifo_U' read by process 'toe_top_toe_top.toe_check_ipv4_checksum_32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_checksumValidFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    36: begin
                        if (~processPseudoHeader_512_U0.rxEng_dataBuffer3a_blk_n) begin
                            if (~rxEng_dataBuffer3a_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer3a_U' written by process 'toe_top_toe_top.rshiftWordByOctet_net_axis_512_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3a_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer3a_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer3a_U' read by process 'toe_top_toe_top.rshiftWordByOctet_net_axis_512_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3a_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    39: begin
                        if (~processPseudoHeader_512_U0.rxEng_headerMetaFifo_blk_n) begin
                            if (~rxEng_headerMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_headerMetaFifo_U' written by process 'toe_top_toe_top.merge_header_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_headerMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_headerMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_headerMetaFifo_U' read by process 'toe_top_toe_top.merge_header_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_headerMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    19: begin
                        if (~processPseudoHeader_512_U0.rxEng2portTable_check_req_blk_n) begin
                            if (~rxEng2portTable_check_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2portTable_check_req_U' written by process 'toe_top_toe_top.check_in_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2portTable_check_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2portTable_check_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2portTable_check_req_U' read by process 'toe_top_toe_top.check_in_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2portTable_check_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    40: begin
                        if (~processPseudoHeader_512_U0.rxEng_tupleBuffer_blk_n) begin
                            if (~rxEng_tupleBuffer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_tupleBuffer_U' written by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_tupleBuffer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_tupleBuffer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_tupleBuffer_U' read by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_tupleBuffer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    37: begin
                        if (~processPseudoHeader_512_U0.rxEng_optionalFieldsMetaFifo_blk_n) begin
                            if (~rxEng_optionalFieldsMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_optionalFieldsMetaFifo_U' written by process 'toe_top_toe_top.drop_optional_header_fields_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_optionalFieldsMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_optionalFieldsMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_optionalFieldsMetaFifo_U' read by process 'toe_top_toe_top.drop_optional_header_fields_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_optionalFieldsMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                36 : begin
                    case(index2)
                    35: begin
                        if (~rshiftWordByOctet_net_axis_512_512_3_U0.rxEng_dataBuffer3a_blk_n) begin
                            if (~rxEng_dataBuffer3a_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer3a_U' written by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3a_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer3a_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer3a_U' read by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3a_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    37: begin
                        if (~rshiftWordByOctet_net_axis_512_512_3_U0.rxEng_dataBuffer3b_blk_n) begin
                            if (~rxEng_dataBuffer3b_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer3b_U' written by process 'toe_top_toe_top.drop_optional_header_fields_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3b_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer3b_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer3b_U' read by process 'toe_top_toe_top.drop_optional_header_fields_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3b_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                37 : begin
                    case(index2)
                    35: begin
                        if (~drop_optional_header_fields_512_U0.rxEng_optionalFieldsMetaFifo_blk_n) begin
                            if (~rxEng_optionalFieldsMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_optionalFieldsMetaFifo_U' written by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_optionalFieldsMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_optionalFieldsMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_optionalFieldsMetaFifo_U' read by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_optionalFieldsMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    36: begin
                        if (~drop_optional_header_fields_512_U0.rxEng_dataBuffer3b_blk_n) begin
                            if (~rxEng_dataBuffer3b_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer3b_U' written by process 'toe_top_toe_top.rshiftWordByOctet_net_axis_512_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3b_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer3b_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer3b_U' read by process 'toe_top_toe_top.rshiftWordByOctet_net_axis_512_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3b_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    42: begin
                        if (~drop_optional_header_fields_512_U0.rxEng_dataBuffer3_blk_n) begin
                            if (~rxEng_dataBuffer3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer3_U' written by process 'toe_top_toe_top.rxPackageDropper_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer3_U' read by process 'toe_top_toe_top.rxPackageDropper_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    38: begin
                        if (~drop_optional_header_fields_512_U0.rxEng_dataOffsetFifo_blk_n) begin
                            if (~rxEng_dataOffsetFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataOffsetFifo_U' written by process 'toe_top_toe_top.parse_optional_header_fields_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataOffsetFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataOffsetFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataOffsetFifo_U' read by process 'toe_top_toe_top.parse_optional_header_fields_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataOffsetFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~drop_optional_header_fields_512_U0.rxEng_optionalFieldsFifo_blk_n) begin
                            if (~rxEng_optionalFieldsFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_optionalFieldsFifo_U' written by process 'toe_top_toe_top.parse_optional_header_fields_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_optionalFieldsFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_optionalFieldsFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_optionalFieldsFifo_U' read by process 'toe_top_toe_top.parse_optional_header_fields_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_optionalFieldsFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                38 : begin
                    case(index2)
                    37: begin
                        if (~parse_optional_header_fields_U0.rxEng_dataOffsetFifo_blk_n) begin
                            if (~rxEng_dataOffsetFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataOffsetFifo_U' written by process 'toe_top_toe_top.drop_optional_header_fields_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataOffsetFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataOffsetFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataOffsetFifo_U' read by process 'toe_top_toe_top.drop_optional_header_fields_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataOffsetFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~parse_optional_header_fields_U0.rxEng_optionalFieldsFifo_blk_n) begin
                            if (~rxEng_optionalFieldsFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_optionalFieldsFifo_U' written by process 'toe_top_toe_top.drop_optional_header_fields_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_optionalFieldsFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_optionalFieldsFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_optionalFieldsFifo_U' read by process 'toe_top_toe_top.drop_optional_header_fields_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_optionalFieldsFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    39: begin
                        if (~parse_optional_header_fields_U0.rxEng_winScaleFifo_blk_n) begin
                            if (~rxEng_winScaleFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_winScaleFifo_U' written by process 'toe_top_toe_top.merge_header_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_winScaleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_winScaleFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_winScaleFifo_U' read by process 'toe_top_toe_top.merge_header_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_winScaleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                39 : begin
                    case(index2)
                    35: begin
                        if (~merge_header_meta_U0.rxEng_headerMetaFifo_blk_n) begin
                            if (~rxEng_headerMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_headerMetaFifo_U' written by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_headerMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_headerMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_headerMetaFifo_U' read by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_headerMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    40: begin
                        if (~merge_header_meta_U0.rxEng_metaDataFifo_blk_n) begin
                            if (~rxEng_metaDataFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_metaDataFifo_U' written by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaDataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_metaDataFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_metaDataFifo_U' read by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaDataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    38: begin
                        if (~merge_header_meta_U0.rxEng_winScaleFifo_blk_n) begin
                            if (~rxEng_winScaleFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_winScaleFifo_U' written by process 'toe_top_toe_top.parse_optional_header_fields_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_winScaleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_winScaleFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_winScaleFifo_U' read by process 'toe_top_toe_top.parse_optional_header_fields_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_winScaleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                40 : begin
                    case(index2)
                    39: begin
                        if (~rxMetadataHandler_U0.rxEng_metaDataFifo_blk_n) begin
                            if (~rxEng_metaDataFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_metaDataFifo_U' written by process 'toe_top_toe_top.merge_header_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaDataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_metaDataFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_metaDataFifo_U' read by process 'toe_top_toe_top.merge_header_meta_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaDataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    20: begin
                        if (~rxMetadataHandler_U0.portTable2rxEng_check_rsp_blk_n) begin
                            if (~portTable2rxEng_check_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.portTable2rxEng_check_rsp_U' written by process 'toe_top_toe_top.check_out_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2rxEng_check_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~portTable2rxEng_check_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.portTable2rxEng_check_rsp_U' read by process 'toe_top_toe_top.check_out_multiplexer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2rxEng_check_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    35: begin
                        if (~rxMetadataHandler_U0.rxEng_tupleBuffer_blk_n) begin
                            if (~rxEng_tupleBuffer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_tupleBuffer_U' written by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_tupleBuffer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_tupleBuffer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_tupleBuffer_U' read by process 'toe_top_toe_top.processPseudoHeader_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_tupleBuffer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    43: begin
                        if (~rxMetadataHandler_U0.rxEng_metaHandlerEventFifo_blk_n) begin
                            if (~rxEng_metaHandlerEventFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_metaHandlerEventFifo_U' written by process 'toe_top_toe_top.rxEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaHandlerEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_metaHandlerEventFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_metaHandlerEventFifo_U' read by process 'toe_top_toe_top.rxEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaHandlerEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    42: begin
                        if (~rxMetadataHandler_U0.rxEng_metaHandlerDropFifo_blk_n) begin
                            if (~rxEng_metaHandlerDropFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_metaHandlerDropFifo_U' written by process 'toe_top_toe_top.rxPackageDropper_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaHandlerDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_metaHandlerDropFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_metaHandlerDropFifo_U' read by process 'toe_top_toe_top.rxPackageDropper_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaHandlerDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    9: begin
                        if (~rxMetadataHandler_U0.rxEng2sLookup_req_blk_n) begin
                            if (~rxEng2sLookup_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2sLookup_req_U' written by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2sLookup_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2sLookup_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2sLookup_req_U' read by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2sLookup_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rxMetadataHandler_U0.sLookup2rxEng_rsp_blk_n) begin
                            if (~sLookup2rxEng_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sLookup2rxEng_rsp_U' written by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2rxEng_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sLookup2rxEng_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sLookup2rxEng_rsp_U' read by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2rxEng_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    41: begin
                        if (~rxMetadataHandler_U0.rxEng_fsmMetaDataFifo_blk_n) begin
                            if (~rxEng_fsmMetaDataFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_fsmMetaDataFifo_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmMetaDataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_fsmMetaDataFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_fsmMetaDataFifo_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmMetaDataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                41 : begin
                    case(index2)
                    0: begin
                        if (~rxTcpFSM_U0.rxbuffer_data_count_blk_n) begin
                            if (~axis_data_count_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.axis_data_count_c_U' written by process 'toe_top_toe_top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.axis_data_count_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~axis_data_count_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.axis_data_count_c_U' read by process 'toe_top_toe_top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.axis_data_count_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rxTcpFSM_U0.rxbuffer_max_data_count_blk_n) begin
                            if (~axis_max_data_count_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.axis_max_data_count_c_U' written by process 'toe_top_toe_top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.axis_max_data_count_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~axis_max_data_count_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.axis_max_data_count_c_U' read by process 'toe_top_toe_top.entry_proc_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.axis_max_data_count_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    40: begin
                        if (~rxTcpFSM_U0.rxEng_fsmMetaDataFifo_blk_n) begin
                            if (~rxEng_fsmMetaDataFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_fsmMetaDataFifo_U' written by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmMetaDataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_fsmMetaDataFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_fsmMetaDataFifo_U' read by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmMetaDataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~rxTcpFSM_U0.rxEng2stateTable_upd_req_blk_n) begin
                            if (~rxEng2stateTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2stateTable_upd_req_U' written by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2stateTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2stateTable_upd_req_U' read by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rxTcpFSM_U0.stateTable2rxEng_upd_rsp_blk_n) begin
                            if (~stateTable2rxEng_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.stateTable2rxEng_upd_rsp_U' written by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2rxEng_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.stateTable2rxEng_upd_rsp_U' read by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    15: begin
                        if (~rxTcpFSM_U0.rxEng2rxSar_upd_req_blk_n) begin
                            if (~rxEng2rxSar_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2rxSar_upd_req_U' written by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2rxSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2rxSar_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2rxSar_upd_req_U' read by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2rxSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rxTcpFSM_U0.rxSar2rxEng_upd_rsp_blk_n) begin
                            if (~rxSar2rxEng_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxSar2rxEng_upd_rsp_U' written by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxSar2rxEng_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxSar2rxEng_upd_rsp_U' read by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    16: begin
                        if (~rxTcpFSM_U0.rxEng2txSar_upd_req_blk_n) begin
                            if (~rxEng2txSar_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2txSar_upd_req_U' written by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2txSar_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2txSar_upd_req_U' read by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rxTcpFSM_U0.txSar2rxEng_upd_rsp_blk_n) begin
                            if (~txSar2rxEng_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txSar2rxEng_upd_rsp_U' written by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txSar2rxEng_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txSar2rxEng_upd_rsp_U' read by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2rxEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    22: begin
                        if (~rxTcpFSM_U0.rxEng2timer_clearRetransmitTimer_blk_n) begin
                            if (~rxEng2timer_clearRetransmitTimer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2timer_clearRetransmitTimer_U' written by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_clearRetransmitTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2timer_clearRetransmitTimer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2timer_clearRetransmitTimer_U' read by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_clearRetransmitTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    23: begin
                        if (~rxTcpFSM_U0.rxEng2timer_clearProbeTimer_blk_n) begin
                            if (~rxEng2timer_clearProbeTimer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2timer_clearProbeTimer_U' written by process 'toe_top_toe_top.probe_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_clearProbeTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2timer_clearProbeTimer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2timer_clearProbeTimer_U' read by process 'toe_top_toe_top.probe_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_clearProbeTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    61: begin
                        if (~rxTcpFSM_U0.rxEng2rxApp_notification_blk_n) begin
                            if (~rxEng2rxApp_notification_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2rxApp_notification_U' written by process 'toe_top_toe_top.stream_merger_appNotification_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2rxApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2rxApp_notification_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2rxApp_notification_U' read by process 'toe_top_toe_top.stream_merger_appNotification_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2rxApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    42: begin
                        if (~rxTcpFSM_U0.rxEng_fsmDropFifo_blk_n) begin
                            if (~rxEng_fsmDropFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_fsmDropFifo_U' written by process 'toe_top_toe_top.rxPackageDropper_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_fsmDropFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_fsmDropFifo_U' read by process 'toe_top_toe_top.rxPackageDropper_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    43: begin
                        if (~rxTcpFSM_U0.rxEng_fsmEventFifo_blk_n) begin
                            if (~rxEng_fsmEventFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_fsmEventFifo_U' written by process 'toe_top_toe_top.rxEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_fsmEventFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_fsmEventFifo_U' read by process 'toe_top_toe_top.rxEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    24: begin
                        if (~rxTcpFSM_U0.rxEng2timer_setCloseTimer_blk_n) begin
                            if (~rxEng2timer_setCloseTimer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2timer_setCloseTimer_U' written by process 'toe_top_toe_top.close_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_setCloseTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2timer_setCloseTimer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2timer_setCloseTimer_U' read by process 'toe_top_toe_top.close_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2timer_setCloseTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    67: begin
                        if (~rxTcpFSM_U0.conEstablishedFifo_blk_n) begin
                            if (~conEstablishedFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.conEstablishedFifo_U' written by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.conEstablishedFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~conEstablishedFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.conEstablishedFifo_U' read by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.conEstablishedFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                42 : begin
                    case(index2)
                    40: begin
                        if (~rxPackageDropper_512_U0.rxEng_metaHandlerDropFifo_blk_n) begin
                            if (~rxEng_metaHandlerDropFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_metaHandlerDropFifo_U' written by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaHandlerDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_metaHandlerDropFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_metaHandlerDropFifo_U' read by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaHandlerDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    41: begin
                        if (~rxPackageDropper_512_U0.rxEng_fsmDropFifo_blk_n) begin
                            if (~rxEng_fsmDropFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_fsmDropFifo_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_fsmDropFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_fsmDropFifo_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmDropFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    37: begin
                        if (~rxPackageDropper_512_U0.rxEng_dataBuffer3_blk_n) begin
                            if (~rxEng_dataBuffer3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_dataBuffer3_U' written by process 'toe_top_toe_top.drop_optional_header_fields_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_dataBuffer3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_dataBuffer3_U' read by process 'toe_top_toe_top.drop_optional_header_fields_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_dataBuffer3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    5: begin
                        if (~rxPackageDropper_512_U0.rxBufferWriteData_internal_blk_n) begin
                            if (~rxBufferWriteData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxBufferWriteData_internal_U' written by process 'toe_top_toe_top.convert_net_axis_to_axis_512_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferWriteData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxBufferWriteData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxBufferWriteData_internal_U' read by process 'toe_top_toe_top.convert_net_axis_to_axis_512_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferWriteData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                43 : begin
                    case(index2)
                    40: begin
                        if (~rxEventMerger_U0.rxEng_metaHandlerEventFifo_blk_n) begin
                            if (~rxEng_metaHandlerEventFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_metaHandlerEventFifo_U' written by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaHandlerEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_metaHandlerEventFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_metaHandlerEventFifo_U' read by process 'toe_top_toe_top.rxMetadataHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_metaHandlerEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    26: begin
                        if (~rxEventMerger_U0.rxEng2eventEng_setEvent_blk_n) begin
                            if (~rxEng2eventEng_setEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2eventEng_setEvent_U' written by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2eventEng_setEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2eventEng_setEvent_U' read by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    41: begin
                        if (~rxEventMerger_U0.rxEng_fsmEventFifo_blk_n) begin
                            if (~rxEng_fsmEventFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng_fsmEventFifo_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng_fsmEventFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng_fsmEventFifo_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng_fsmEventFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                44 : begin
                    case(index2)
                    27: begin
                        if (~metaLoader_U0.eventEng2txEng_event_blk_n) begin
                            if (~eventEng2txEng_event_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.eventEng2txEng_event_U' written by process 'toe_top_toe_top.ack_delay_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.eventEng2txEng_event_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~eventEng2txEng_event_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.eventEng2txEng_event_U' read by process 'toe_top_toe_top.ack_delay_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.eventEng2txEng_event_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    26: begin
                        if (~metaLoader_U0.txEngFifoReadCount_blk_n) begin
                            if (~txEngFifoReadCount_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEngFifoReadCount_U' written by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEngFifoReadCount_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEngFifoReadCount_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEngFifoReadCount_U' read by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEngFifoReadCount_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    15: begin
                        if (~metaLoader_U0.txEng2rxSar_req_blk_n) begin
                            if (~txEng2rxSar_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng2rxSar_req_U' written by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2rxSar_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng2rxSar_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng2rxSar_req_U' read by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2rxSar_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~metaLoader_U0.rxSar2txEng_rsp_blk_n) begin
                            if (~rxSar2txEng_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxSar2txEng_rsp_U' written by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2txEng_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxSar2txEng_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxSar2txEng_rsp_U' read by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2txEng_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    16: begin
                        if (~metaLoader_U0.txEng2txSar_upd_req_blk_n) begin
                            if (~txEng2txSar_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng2txSar_upd_req_U' written by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng2txSar_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng2txSar_upd_req_U' read by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~metaLoader_U0.txSar2txEng_upd_rsp_blk_n) begin
                            if (~txSar2txEng_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txSar2txEng_upd_rsp_U' written by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txSar2txEng_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txSar2txEng_upd_rsp_U' read by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txEng_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    23: begin
                        if (~metaLoader_U0.txEng2timer_setProbeTimer_blk_n) begin
                            if (~txEng2timer_setProbeTimer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng2timer_setProbeTimer_U' written by process 'toe_top_toe_top.probe_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2timer_setProbeTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng2timer_setProbeTimer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng2timer_setProbeTimer_U' read by process 'toe_top_toe_top.probe_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2timer_setProbeTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    57: begin
                        if (~metaLoader_U0.txEng_ipMetaFifo_blk_n) begin
                            if (~txEng_ipMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_ipMetaFifo_U' written by process 'toe_top_toe_top.generate_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_ipMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_ipMetaFifo_U' read by process 'toe_top_toe_top.generate_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    50: begin
                        if (~metaLoader_U0.txEng_tcpMetaFifo_blk_n) begin
                            if (~txEng_tcpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpMetaFifo_U' written by process 'toe_top_toe_top.pseudoHeaderConstructionNew_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpMetaFifo_U' read by process 'toe_top_toe_top.pseudoHeaderConstructionNew_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    46: begin
                        if (~metaLoader_U0.txEng_isLookUpFifo_blk_n) begin
                            if (~txEng_isLookUpFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_isLookUpFifo_U' written by process 'toe_top_toe_top.tupleSplitter_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_isLookUpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_isLookUpFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_isLookUpFifo_U' read by process 'toe_top_toe_top.tupleSplitter_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_isLookUpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~metaLoader_U0.txEng_tupleShortCutFifo_blk_n) begin
                            if (~txEng_tupleShortCutFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tupleShortCutFifo_U' written by process 'toe_top_toe_top.tupleSplitter_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tupleShortCutFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tupleShortCutFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tupleShortCutFifo_U' read by process 'toe_top_toe_top.tupleSplitter_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tupleShortCutFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    48: begin
                        if (~metaLoader_U0.txEng_isDDRbypass_blk_n) begin
                            if (~txEng_isDDRbypass_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_isDDRbypass_U' written by process 'toe_top_toe_top.read_data_arbiter_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_isDDRbypass_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_isDDRbypass_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_isDDRbypass_U' read by process 'toe_top_toe_top.read_data_arbiter_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_isDDRbypass_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~metaLoader_U0.txEng2sLookup_rev_req_blk_n) begin
                            if (~txEng2sLookup_rev_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng2sLookup_rev_req_U' written by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2sLookup_rev_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng2sLookup_rev_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng2sLookup_rev_req_U' read by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2sLookup_rev_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    22: begin
                        if (~metaLoader_U0.txEng2timer_setRetransmitTimer_blk_n) begin
                            if (~txEng2timer_setRetransmitTimer_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng2timer_setRetransmitTimer_U' written by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2timer_setRetransmitTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng2timer_setRetransmitTimer_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng2timer_setRetransmitTimer_U' read by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng2timer_setRetransmitTimer_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    45: begin
                        if (~metaLoader_U0.txMetaloader2memAccessBreakdown_blk_n) begin
                            if (~txMetaloader2memAccessBreakdown_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txMetaloader2memAccessBreakdown_U' written by process 'toe_top_toe_top.txEngMemAccessBreakdown_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txMetaloader2memAccessBreakdown_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txMetaloader2memAccessBreakdown_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txMetaloader2memAccessBreakdown_U' read by process 'toe_top_toe_top.txEngMemAccessBreakdown_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txMetaloader2memAccessBreakdown_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                45 : begin
                    case(index2)
                    44: begin
                        if (~txEngMemAccessBreakdown_U0.txMetaloader2memAccessBreakdown_blk_n) begin
                            if (~txMetaloader2memAccessBreakdown_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txMetaloader2memAccessBreakdown_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txMetaloader2memAccessBreakdown_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txMetaloader2memAccessBreakdown_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txMetaloader2memAccessBreakdown_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txMetaloader2memAccessBreakdown_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    47: begin
                        if (~txEngMemAccessBreakdown_U0.memAccessBreakdown2txPkgStitcher_blk_n) begin
                            if (~memAccessBreakdown2txPkgStitcher_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.memAccessBreakdown2txPkgStitcher_U' written by process 'toe_top_toe_top.read_data_stitching_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.memAccessBreakdown2txPkgStitcher_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~memAccessBreakdown2txPkgStitcher_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.memAccessBreakdown2txPkgStitcher_U' read by process 'toe_top_toe_top.read_data_stitching_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.memAccessBreakdown2txPkgStitcher_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                46 : begin
                    case(index2)
                    44: begin
                        if (~tupleSplitter_U0.txEng_isLookUpFifo_blk_n) begin
                            if (~txEng_isLookUpFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_isLookUpFifo_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_isLookUpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_isLookUpFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_isLookUpFifo_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_isLookUpFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~tupleSplitter_U0.txEng_tupleShortCutFifo_blk_n) begin
                            if (~txEng_tupleShortCutFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tupleShortCutFifo_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tupleShortCutFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tupleShortCutFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tupleShortCutFifo_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tupleShortCutFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    13: begin
                        if (~tupleSplitter_U0.sLookup2txEng_rev_rsp_blk_n) begin
                            if (~sLookup2txEng_rev_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sLookup2txEng_rev_rsp_U' written by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2txEng_rev_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sLookup2txEng_rev_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sLookup2txEng_rev_rsp_U' read by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2txEng_rev_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    57: begin
                        if (~tupleSplitter_U0.txEng_ipTupleFifo_blk_n) begin
                            if (~txEng_ipTupleFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_ipTupleFifo_U' written by process 'toe_top_toe_top.generate_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_ipTupleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_ipTupleFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_ipTupleFifo_U' read by process 'toe_top_toe_top.generate_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_ipTupleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    50: begin
                        if (~tupleSplitter_U0.txEng_tcpTupleFifo_blk_n) begin
                            if (~txEng_tcpTupleFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpTupleFifo_U' written by process 'toe_top_toe_top.pseudoHeaderConstructionNew_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpTupleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpTupleFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpTupleFifo_U' read by process 'toe_top_toe_top.pseudoHeaderConstructionNew_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpTupleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                47 : begin
                    case(index2)
                    45: begin
                        if (~read_data_stitching_512_U0.memAccessBreakdown2txPkgStitcher_blk_n) begin
                            if (~memAccessBreakdown2txPkgStitcher_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.memAccessBreakdown2txPkgStitcher_U' written by process 'toe_top_toe_top.txEngMemAccessBreakdown_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.memAccessBreakdown2txPkgStitcher_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~memAccessBreakdown2txPkgStitcher_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.memAccessBreakdown2txPkgStitcher_U' read by process 'toe_top_toe_top.txEngMemAccessBreakdown_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.memAccessBreakdown2txPkgStitcher_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    3: begin
                        if (~read_data_stitching_512_U0.txBufferReadData_internal_blk_n) begin
                            if (~txBufferReadData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txBufferReadData_internal_U' written by process 'toe_top_toe_top.convert_axis_to_net_axis_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferReadData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txBufferReadData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txBufferReadData_internal_U' read by process 'toe_top_toe_top.convert_axis_to_net_axis_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferReadData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    48: begin
                        if (~read_data_stitching_512_U0.txBufferReadDataStitched_blk_n) begin
                            if (~txBufferReadDataStitched_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txBufferReadDataStitched_U' written by process 'toe_top_toe_top.read_data_arbiter_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferReadDataStitched_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txBufferReadDataStitched_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txBufferReadDataStitched_U' read by process 'toe_top_toe_top.read_data_arbiter_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferReadDataStitched_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                48 : begin
                    case(index2)
                    44: begin
                        if (~read_data_arbiter_512_U0.txEng_isDDRbypass_blk_n) begin
                            if (~txEng_isDDRbypass_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_isDDRbypass_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_isDDRbypass_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_isDDRbypass_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_isDDRbypass_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_isDDRbypass_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    47: begin
                        if (~read_data_arbiter_512_U0.txBufferReadDataStitched_blk_n) begin
                            if (~txBufferReadDataStitched_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txBufferReadDataStitched_U' written by process 'toe_top_toe_top.read_data_stitching_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferReadDataStitched_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txBufferReadDataStitched_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txBufferReadDataStitched_U' read by process 'toe_top_toe_top.read_data_stitching_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferReadDataStitched_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    49: begin
                        if (~read_data_arbiter_512_U0.txEng_tcpPkgBuffer0_blk_n) begin
                            if (~txEng_tcpPkgBuffer0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer0_U' written by process 'toe_top_toe_top.lshiftWordByOctet_512_51_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer0_U' read by process 'toe_top_toe_top.lshiftWordByOctet_512_51_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    65: begin
                        if (~read_data_arbiter_512_U0.txApp2txEng_data_stream_blk_n) begin
                            if (~txApp2txEng_data_stream_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2txEng_data_stream_U' written by process 'toe_top_toe_top.toe_duplicate_stream_net_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txEng_data_stream_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2txEng_data_stream_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2txEng_data_stream_U' read by process 'toe_top_toe_top.toe_duplicate_stream_net_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txEng_data_stream_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                49 : begin
                    case(index2)
                    50: begin
                        if (~lshiftWordByOctet_512_51_U0.txEng_shift2pseudoFifo_blk_n) begin
                            if (~txEng_shift2pseudoFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_shift2pseudoFifo_U' written by process 'toe_top_toe_top.pseudoHeaderConstructionNew_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_shift2pseudoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_shift2pseudoFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_shift2pseudoFifo_U' read by process 'toe_top_toe_top.pseudoHeaderConstructionNew_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_shift2pseudoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    48: begin
                        if (~lshiftWordByOctet_512_51_U0.txEng_tcpPkgBuffer0_blk_n) begin
                            if (~txEng_tcpPkgBuffer0_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer0_U' written by process 'toe_top_toe_top.read_data_arbiter_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer0_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer0_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer0_U' read by process 'toe_top_toe_top.read_data_arbiter_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer0_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                50 : begin
                    case(index2)
                    44: begin
                        if (~pseudoHeaderConstructionNew_512_U0.txEng_tcpMetaFifo_blk_n) begin
                            if (~txEng_tcpMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpMetaFifo_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpMetaFifo_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    46: begin
                        if (~pseudoHeaderConstructionNew_512_U0.txEng_tcpTupleFifo_blk_n) begin
                            if (~txEng_tcpTupleFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpTupleFifo_U' written by process 'toe_top_toe_top.tupleSplitter_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpTupleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpTupleFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpTupleFifo_U' read by process 'toe_top_toe_top.tupleSplitter_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpTupleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    51: begin
                        if (~pseudoHeaderConstructionNew_512_U0.txEng_tcpPkgBuffer1_blk_n) begin
                            if (~txEng_tcpPkgBuffer1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer1_U' written by process 'toe_top_toe_top.two_complement_subchecksums_512_22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer1_U' read by process 'toe_top_toe_top.two_complement_subchecksums_512_22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    49: begin
                        if (~pseudoHeaderConstructionNew_512_U0.txEng_shift2pseudoFifo_blk_n) begin
                            if (~txEng_shift2pseudoFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_shift2pseudoFifo_U' written by process 'toe_top_toe_top.lshiftWordByOctet_512_51_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_shift2pseudoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_shift2pseudoFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_shift2pseudoFifo_U' read by process 'toe_top_toe_top.lshiftWordByOctet_512_51_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_shift2pseudoFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                51 : begin
                    case(index2)
                    50: begin
                        if (~two_complement_subchecksums_512_22_U0.txEng_tcpPkgBuffer1_blk_n) begin
                            if (~txEng_tcpPkgBuffer1_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer1_U' written by process 'toe_top_toe_top.pseudoHeaderConstructionNew_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer1_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer1_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer1_U' read by process 'toe_top_toe_top.pseudoHeaderConstructionNew_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer1_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    53: begin
                        if (~two_complement_subchecksums_512_22_U0.txEng_tcpPkgBuffer2_blk_n) begin
                            if (~txEng_tcpPkgBuffer2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer2_U' written by process 'toe_top_toe_top.remove_pseudo_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer2_U' read by process 'toe_top_toe_top.remove_pseudo_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    52: begin
                        if (~two_complement_subchecksums_512_22_U0.txEng_subChecksumsFifo_blk_n) begin
                            if (~txEng_subChecksumsFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_subChecksumsFifo_U' written by process 'toe_top_toe_top.finalize_ipv4_checksum_32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_subChecksumsFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_subChecksumsFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_subChecksumsFifo_U' read by process 'toe_top_toe_top.finalize_ipv4_checksum_32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_subChecksumsFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                52 : begin
                    case(index2)
                    51: begin
                        if (~finalize_ipv4_checksum_32_U0.txEng_subChecksumsFifo_blk_n) begin
                            if (~txEng_subChecksumsFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_subChecksumsFifo_U' written by process 'toe_top_toe_top.two_complement_subchecksums_512_22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_subChecksumsFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_subChecksumsFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_subChecksumsFifo_U' read by process 'toe_top_toe_top.two_complement_subchecksums_512_22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_subChecksumsFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    55: begin
                        if (~finalize_ipv4_checksum_32_U0.txEng_tcpChecksumFifo_blk_n) begin
                            if (~txEng_tcpChecksumFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpChecksumFifo_U' written by process 'toe_top_toe_top.insert_checksum_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpChecksumFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpChecksumFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpChecksumFifo_U' read by process 'toe_top_toe_top.insert_checksum_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpChecksumFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                53 : begin
                    case(index2)
                    51: begin
                        if (~remove_pseudo_header_512_U0.txEng_tcpPkgBuffer2_blk_n) begin
                            if (~txEng_tcpPkgBuffer2_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer2_U' written by process 'toe_top_toe_top.two_complement_subchecksums_512_22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer2_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer2_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer2_U' read by process 'toe_top_toe_top.two_complement_subchecksums_512_22_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer2_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    54: begin
                        if (~remove_pseudo_header_512_U0.txEng_tcpPkgBuffer3_blk_n) begin
                            if (~txEng_tcpPkgBuffer3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer3_U' written by process 'toe_top_toe_top.rshiftWordByOctet_net_axis_512_512_53_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer3_U' read by process 'toe_top_toe_top.rshiftWordByOctet_net_axis_512_512_53_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                54 : begin
                    case(index2)
                    53: begin
                        if (~rshiftWordByOctet_net_axis_512_512_53_U0.txEng_tcpPkgBuffer3_blk_n) begin
                            if (~txEng_tcpPkgBuffer3_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer3_U' written by process 'toe_top_toe_top.remove_pseudo_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer3_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer3_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer3_U' read by process 'toe_top_toe_top.remove_pseudo_header_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer3_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    55: begin
                        if (~rshiftWordByOctet_net_axis_512_512_53_U0.txEng_tcpPkgBuffer4_blk_n) begin
                            if (~txEng_tcpPkgBuffer4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer4_U' written by process 'toe_top_toe_top.insert_checksum_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer4_U' read by process 'toe_top_toe_top.insert_checksum_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                55 : begin
                    case(index2)
                    52: begin
                        if (~insert_checksum_512_U0.txEng_tcpChecksumFifo_blk_n) begin
                            if (~txEng_tcpChecksumFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpChecksumFifo_U' written by process 'toe_top_toe_top.finalize_ipv4_checksum_32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpChecksumFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpChecksumFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpChecksumFifo_U' read by process 'toe_top_toe_top.finalize_ipv4_checksum_32_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpChecksumFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    54: begin
                        if (~insert_checksum_512_U0.txEng_tcpPkgBuffer4_blk_n) begin
                            if (~txEng_tcpPkgBuffer4_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer4_U' written by process 'toe_top_toe_top.rshiftWordByOctet_net_axis_512_512_53_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer4_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer4_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer4_U' read by process 'toe_top_toe_top.rshiftWordByOctet_net_axis_512_512_53_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer4_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    56: begin
                        if (~insert_checksum_512_U0.txEng_tcpPkgBuffer5_blk_n) begin
                            if (~txEng_tcpPkgBuffer5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer5_U' written by process 'toe_top_toe_top.lshiftWordByOctet_512_52_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer5_U' read by process 'toe_top_toe_top.lshiftWordByOctet_512_52_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                56 : begin
                    case(index2)
                    57: begin
                        if (~lshiftWordByOctet_512_52_U0.txEng_tcpPkgBuffer6_blk_n) begin
                            if (~txEng_tcpPkgBuffer6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer6_U' written by process 'toe_top_toe_top.generate_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer6_U' read by process 'toe_top_toe_top.generate_ipv4_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    55: begin
                        if (~lshiftWordByOctet_512_52_U0.txEng_tcpPkgBuffer5_blk_n) begin
                            if (~txEng_tcpPkgBuffer5_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer5_U' written by process 'toe_top_toe_top.insert_checksum_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer5_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer5_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer5_U' read by process 'toe_top_toe_top.insert_checksum_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer5_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                57 : begin
                    case(index2)
                    44: begin
                        if (~generate_ipv4_512_U0.txEng_ipMetaFifo_blk_n) begin
                            if (~txEng_ipMetaFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_ipMetaFifo_U' written by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_ipMetaFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_ipMetaFifo_U' read by process 'toe_top_toe_top.metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_ipMetaFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    46: begin
                        if (~generate_ipv4_512_U0.txEng_ipTupleFifo_blk_n) begin
                            if (~txEng_ipTupleFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_ipTupleFifo_U' written by process 'toe_top_toe_top.tupleSplitter_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_ipTupleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_ipTupleFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_ipTupleFifo_U' read by process 'toe_top_toe_top.tupleSplitter_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_ipTupleFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    4: begin
                        if (~generate_ipv4_512_U0.ipTxData_internal_blk_n) begin
                            if (~ipTxData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.ipTxData_internal_U' written by process 'toe_top_toe_top.convert_net_axis_to_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ipTxData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~ipTxData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.ipTxData_internal_U' read by process 'toe_top_toe_top.convert_net_axis_to_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.ipTxData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    56: begin
                        if (~generate_ipv4_512_U0.txEng_tcpPkgBuffer6_blk_n) begin
                            if (~txEng_tcpPkgBuffer6_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer6_U' written by process 'toe_top_toe_top.lshiftWordByOctet_512_52_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer6_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txEng_tcpPkgBuffer6_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txEng_tcpPkgBuffer6_U' read by process 'toe_top_toe_top.lshiftWordByOctet_512_52_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txEng_tcpPkgBuffer6_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                58 : begin
                    case(index2)
                    15: begin
                        if (~rx_app_stream_if_U0.rxApp2rxSar_upd_req_blk_n) begin
                            if (~rxApp2rxSar_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxApp2rxSar_upd_req_U' written by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxApp2rxSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxApp2rxSar_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxApp2rxSar_upd_req_U' read by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxApp2rxSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rx_app_stream_if_U0.rxSar2rxApp_upd_rsp_blk_n) begin
                            if (~rxSar2rxApp_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxSar2rxApp_upd_rsp_U' written by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2rxApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxSar2rxApp_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxSar2rxApp_upd_rsp_U' read by process 'toe_top_toe_top.rx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxSar2rxApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    59: begin
                        if (~rx_app_stream_if_U0.rxBufferReadCmd_blk_n) begin
                            if (~rxBufferReadCmd_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxBufferReadCmd_U' written by process 'toe_top_toe_top.rxAppMemDataRead_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferReadCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxBufferReadCmd_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxBufferReadCmd_U' read by process 'toe_top_toe_top.rxAppMemDataRead_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferReadCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                59 : begin
                    case(index2)
                    58: begin
                        if (~rxAppMemDataRead_512_U0.rxBufferReadCmd_blk_n) begin
                            if (~rxBufferReadCmd_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxBufferReadCmd_U' written by process 'toe_top_toe_top.rx_app_stream_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferReadCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxBufferReadCmd_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxBufferReadCmd_U' read by process 'toe_top_toe_top.rx_app_stream_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferReadCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    2: begin
                        if (~rxAppMemDataRead_512_U0.rxBufferReadData_internal_blk_n) begin
                            if (~rxBufferReadData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxBufferReadData_internal_U' written by process 'toe_top_toe_top.convert_axis_to_net_axis_512_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferReadData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxBufferReadData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxBufferReadData_internal_U' read by process 'toe_top_toe_top.convert_axis_to_net_axis_512_1_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxBufferReadData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    8: begin
                        if (~rxAppMemDataRead_512_U0.rxDataRsp_internal_blk_n) begin
                            if (~rxDataRsp_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxDataRsp_internal_U' written by process 'toe_top_toe_top.convert_net_axis_to_axis_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxDataRsp_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxDataRsp_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxDataRsp_internal_U' read by process 'toe_top_toe_top.convert_net_axis_to_axis_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxDataRsp_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                60 : begin
                    case(index2)
                    17: begin
                        if (~rx_app_if_U0.rxApp2portTable_listen_req_blk_n) begin
                            if (~rxApp2portTable_listen_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxApp2portTable_listen_req_U' written by process 'toe_top_toe_top.listening_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxApp2portTable_listen_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxApp2portTable_listen_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxApp2portTable_listen_req_U' read by process 'toe_top_toe_top.listening_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxApp2portTable_listen_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~rx_app_if_U0.portTable2rxApp_listen_rsp_blk_n) begin
                            if (~portTable2rxApp_listen_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.portTable2rxApp_listen_rsp_U' written by process 'toe_top_toe_top.listening_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2rxApp_listen_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~portTable2rxApp_listen_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.portTable2rxApp_listen_rsp_U' read by process 'toe_top_toe_top.listening_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2rxApp_listen_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                61 : begin
                    case(index2)
                    41: begin
                        if (~stream_merger_appNotification_U0.rxEng2rxApp_notification_blk_n) begin
                            if (~rxEng2rxApp_notification_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.rxEng2rxApp_notification_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2rxApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~rxEng2rxApp_notification_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.rxEng2rxApp_notification_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.rxEng2rxApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    22: begin
                        if (~stream_merger_appNotification_U0.timer2rxApp_notification_blk_n) begin
                            if (~timer2rxApp_notification_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.timer2rxApp_notification_U' written by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2rxApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~timer2rxApp_notification_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.timer2rxApp_notification_U' read by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2rxApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                62 : begin
                    case(index2)
                    67: begin
                        if (~txEventMerger_U0.txApp2eventEng_mergeEvent_blk_n) begin
                            if (~txApp2eventEng_mergeEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2eventEng_mergeEvent_U' written by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2eventEng_mergeEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2eventEng_mergeEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2eventEng_mergeEvent_U' read by process 'toe_top_toe_top.tx_app_if_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2eventEng_mergeEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    26: begin
                        if (~txEventMerger_U0.txApp2eventEng_setEvent_blk_n) begin
                            if (~txApp2eventEng_setEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2eventEng_setEvent_U' written by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2eventEng_setEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2eventEng_setEvent_U' read by process 'toe_top_toe_top.event_engine_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2eventEng_setEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    64: begin
                        if (~txEventMerger_U0.txAppStream2event_mergeEvent_blk_n) begin
                            if (~txAppStream2event_mergeEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txAppStream2event_mergeEvent_U' written by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txAppStream2event_mergeEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txAppStream2event_mergeEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txAppStream2event_mergeEvent_U' read by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txAppStream2event_mergeEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    63: begin
                        if (~txEventMerger_U0.txApp_txEventCache_blk_n) begin
                            if (~txApp_txEventCache_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp_txEventCache_U' written by process 'toe_top_toe_top.txAppStatusHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp_txEventCache_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp_txEventCache_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp_txEventCache_U' read by process 'toe_top_toe_top.txAppStatusHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp_txEventCache_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                63 : begin
                    case(index2)
                    62: begin
                        if (~txAppStatusHandler_U0.txApp_txEventCache_blk_n) begin
                            if (~txApp_txEventCache_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp_txEventCache_U' written by process 'toe_top_toe_top.txEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp_txEventCache_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp_txEventCache_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp_txEventCache_U' read by process 'toe_top_toe_top.txEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp_txEventCache_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    16: begin
                        if (~txAppStatusHandler_U0.txApp2txSar_push_blk_n) begin
                            if (~txApp2txSar_push_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2txSar_push_U' written by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txSar_push_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2txSar_push_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2txSar_push_U' read by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txSar_push_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                64 : begin
                    case(index2)
                    14: begin
                        if (~tasi_metaLoader_U0.txApp2stateTable_req_blk_n) begin
                            if (~txApp2stateTable_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2stateTable_req_U' written by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2stateTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2stateTable_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2stateTable_req_U' read by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2stateTable_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~tasi_metaLoader_U0.stateTable2txApp_rsp_blk_n) begin
                            if (~stateTable2txApp_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.stateTable2txApp_rsp_U' written by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2txApp_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2txApp_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.stateTable2txApp_rsp_U' read by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2txApp_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    68: begin
                        if (~tasi_metaLoader_U0.txApp2txSar_upd_req_blk_n) begin
                            if (~txApp2txSar_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2txSar_upd_req_U' written by process 'toe_top_toe_top.tx_app_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2txSar_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2txSar_upd_req_U' read by process 'toe_top_toe_top.tx_app_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~tasi_metaLoader_U0.txSar2txApp_upd_rsp_blk_n) begin
                            if (~txSar2txApp_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txSar2txApp_upd_rsp_U' written by process 'toe_top_toe_top.tx_app_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txSar2txApp_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txSar2txApp_upd_rsp_U' read by process 'toe_top_toe_top.tx_app_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    66: begin
                        if (~tasi_metaLoader_U0.tasi_meta2pkgPushCmd_blk_n) begin
                            if (~tasi_meta2pkgPushCmd_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.tasi_meta2pkgPushCmd_U' written by process 'toe_top_toe_top.tasi_pkg_pusher_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.tasi_meta2pkgPushCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tasi_meta2pkgPushCmd_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.tasi_meta2pkgPushCmd_U' read by process 'toe_top_toe_top.tasi_pkg_pusher_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.tasi_meta2pkgPushCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    62: begin
                        if (~tasi_metaLoader_U0.txAppStream2event_mergeEvent_blk_n) begin
                            if (~txAppStream2event_mergeEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txAppStream2event_mergeEvent_U' written by process 'toe_top_toe_top.txEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txAppStream2event_mergeEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txAppStream2event_mergeEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txAppStream2event_mergeEvent_U' read by process 'toe_top_toe_top.txEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txAppStream2event_mergeEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                65 : begin
                    case(index2)
                    7: begin
                        if (~toe_duplicate_stream_net_axis_512_U0.txDataReq_internal_blk_n) begin
                            if (~txDataReq_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txDataReq_internal_U' written by process 'toe_top_toe_top.convert_axis_to_net_axis_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txDataReq_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txDataReq_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txDataReq_internal_U' read by process 'toe_top_toe_top.convert_axis_to_net_axis_512_3_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txDataReq_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    66: begin
                        if (~toe_duplicate_stream_net_axis_512_U0.tasi_dataFifo_blk_n) begin
                            if (~tasi_dataFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.tasi_dataFifo_U' written by process 'toe_top_toe_top.tasi_pkg_pusher_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.tasi_dataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tasi_dataFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.tasi_dataFifo_U' read by process 'toe_top_toe_top.tasi_pkg_pusher_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.tasi_dataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    48: begin
                        if (~toe_duplicate_stream_net_axis_512_U0.txApp2txEng_data_stream_blk_n) begin
                            if (~txApp2txEng_data_stream_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2txEng_data_stream_U' written by process 'toe_top_toe_top.read_data_arbiter_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txEng_data_stream_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2txEng_data_stream_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2txEng_data_stream_U' read by process 'toe_top_toe_top.read_data_arbiter_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txEng_data_stream_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                66 : begin
                    case(index2)
                    64: begin
                        if (~tasi_pkg_pusher_512_U0.tasi_meta2pkgPushCmd_blk_n) begin
                            if (~tasi_meta2pkgPushCmd_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.tasi_meta2pkgPushCmd_U' written by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.tasi_meta2pkgPushCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tasi_meta2pkgPushCmd_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.tasi_meta2pkgPushCmd_U' read by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.tasi_meta2pkgPushCmd_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    65: begin
                        if (~tasi_pkg_pusher_512_U0.tasi_dataFifo_blk_n) begin
                            if (~tasi_dataFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.tasi_dataFifo_U' written by process 'toe_top_toe_top.toe_duplicate_stream_net_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.tasi_dataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~tasi_dataFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.tasi_dataFifo_U' read by process 'toe_top_toe_top.toe_duplicate_stream_net_axis_512_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.tasi_dataFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    6: begin
                        if (~tasi_pkg_pusher_512_U0.txBufferWriteData_internal_blk_n) begin
                            if (~txBufferWriteData_internal_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txBufferWriteData_internal_U' written by process 'toe_top_toe_top.convert_net_axis_to_axis_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferWriteData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txBufferWriteData_internal_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txBufferWriteData_internal_U' read by process 'toe_top_toe_top.convert_net_axis_to_axis_512_2_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txBufferWriteData_internal_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                67 : begin
                    case(index2)
                    13: begin
                        if (~tx_app_if_U0.myIpAddress_blk_n) begin
                            if (~myIpAddress_c_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.myIpAddress_c_U' written by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.myIpAddress_c_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~myIpAddress_c_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.myIpAddress_c_U' read by process 'toe_top_toe_top.reverseLookupTableInterface_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.myIpAddress_c_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    18: begin
                        if (~tx_app_if_U0.portTable2txApp_port_rsp_blk_n) begin
                            if (~portTable2txApp_port_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.portTable2txApp_port_rsp_U' written by process 'toe_top_toe_top.free_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2txApp_port_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~portTable2txApp_port_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.portTable2txApp_port_rsp_U' read by process 'toe_top_toe_top.free_port_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.portTable2txApp_port_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    9: begin
                        if (~tx_app_if_U0.txApp2sLookup_req_blk_n) begin
                            if (~txApp2sLookup_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2sLookup_req_U' written by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2sLookup_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2sLookup_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2sLookup_req_U' read by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2sLookup_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~tx_app_if_U0.sLookup2txApp_rsp_blk_n) begin
                            if (~sLookup2txApp_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.sLookup2txApp_rsp_U' written by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2txApp_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~sLookup2txApp_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.sLookup2txApp_rsp_U' read by process 'toe_top_toe_top.lookupReplyHandler_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.sLookup2txApp_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    62: begin
                        if (~tx_app_if_U0.txApp2eventEng_mergeEvent_blk_n) begin
                            if (~txApp2eventEng_mergeEvent_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2eventEng_mergeEvent_U' written by process 'toe_top_toe_top.txEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2eventEng_mergeEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2eventEng_mergeEvent_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2eventEng_mergeEvent_U' read by process 'toe_top_toe_top.txEventMerger_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2eventEng_mergeEvent_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    14: begin
                        if (~tx_app_if_U0.txApp2stateTable_upd_req_blk_n) begin
                            if (~txApp2stateTable_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2stateTable_upd_req_U' written by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2stateTable_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2stateTable_upd_req_U' read by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2stateTable_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~tx_app_if_U0.stateTable2txApp_upd_rsp_blk_n) begin
                            if (~stateTable2txApp_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.stateTable2txApp_upd_rsp_U' written by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2txApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~stateTable2txApp_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.stateTable2txApp_upd_rsp_U' read by process 'toe_top_toe_top.state_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.stateTable2txApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    41: begin
                        if (~tx_app_if_U0.conEstablishedFifo_blk_n) begin
                            if (~conEstablishedFifo_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.conEstablishedFifo_U' written by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.conEstablishedFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~conEstablishedFifo_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.conEstablishedFifo_U' read by process 'toe_top_toe_top.rxTcpFSM_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.conEstablishedFifo_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    22: begin
                        if (~tx_app_if_U0.timer2txApp_notification_blk_n) begin
                            if (~timer2txApp_notification_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.timer2txApp_notification_U' written by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2txApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~timer2txApp_notification_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.timer2txApp_notification_U' read by process 'toe_top_toe_top.retransmit_timer_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.timer2txApp_notification_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
                68 : begin
                    case(index2)
                    16: begin
                        if (~tx_app_table_U0.txSar2txApp_ack_push_blk_n) begin
                            if (~txSar2txApp_ack_push_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txSar2txApp_ack_push_U' written by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txApp_ack_push_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txSar2txApp_ack_push_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txSar2txApp_ack_push_U' read by process 'toe_top_toe_top.tx_sar_table_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txApp_ack_push_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    64: begin
                        if (~tx_app_table_U0.txApp2txSar_upd_req_blk_n) begin
                            if (~txApp2txSar_upd_req_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txApp2txSar_upd_req_U' written by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txApp2txSar_upd_req_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txApp2txSar_upd_req_U' read by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txApp2txSar_upd_req_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                        if (~tx_app_table_U0.txSar2txApp_upd_rsp_blk_n) begin
                            if (~txSar2txApp_upd_rsp_U.if_empty_n) begin
                                $display("//      Blocked by empty input FIFO 'toe_top_toe_top.txSar2txApp_upd_rsp_U' written by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status EMPTY");
                            end
                            else if (~txSar2txApp_upd_rsp_U.if_full_n) begin
                                $display("//      Blocked by full output FIFO 'toe_top_toe_top.txSar2txApp_upd_rsp_U' read by process 'toe_top_toe_top.tasi_metaLoader_U0'");
                                $fdisplay(fp, "Dependence_Channel_path toe_top_toe_top.txSar2txApp_upd_rsp_U");
                                $fdisplay(fp, "Dependence_Channel_status FULL");
                            end
                        end
                    end
                    endcase
                end
            endcase
        end
    endtask

    // report
    initial begin : report_deadlock
        integer cycle_id;
        integer cycle_comp_id;
        integer record_time;
        wait (dl_reset == 1);
        cycle_id = 1;
        record_time = 0;
        while (1) begin
            @ (negedge dl_clock);
            case (CS_fsm)
                ST_DL_DETECTED: begin
                    cycle_comp_id = 2;
                    if (dl_detect_reg != dl_done_reg) begin
                        if (dl_done_reg == 'b0) begin
                            print_dl_head;
                            record_time = $time;
                        end
                        print_cycle_start(proc_path(origin), cycle_id);
                        cycle_id = cycle_id + 1;
                    end
                    else begin
                        print_dl_end((cycle_id - 1),record_time);
                        @(negedge dl_clock);
                        @(negedge dl_clock);
                        $finish;
                    end
                end
                ST_DL_REPORT: begin
                    if ((|(dl_in_vec)) & ~(|(dl_in_vec & origin_reg))) begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                        print_cycle_proc_comp(proc_path(dl_in_vec), cycle_comp_id);
                        cycle_comp_id = cycle_comp_id + 1;
                    end
                    else begin
                        print_cycle_chan_comp(dl_in_vec_reg, dl_in_vec);
                    end
                end
            endcase
        end
    end
 
